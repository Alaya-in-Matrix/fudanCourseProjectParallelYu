
module top ( clk, reset, ins_code2_proc2, ins_code1_proc1, pc_proc1_code1, 
        pc_proc2_code2 );
  input [23:0] ins_code2_proc2;
  input [23:0] ins_code1_proc1;
  output [7:0] pc_proc1_code1;
  output [7:0] pc_proc2_code2;
  input clk, reset;
  wire   en_C1_P1, en_C2_P2, en_M_C1, msg_C2_C1, allowRead_C2_C1, rm_C2_C1,
         wm_C2_C1, msg_C1_C2, allowRead_C1_C2, rm_C1_C2, wm_C1_C2, en_M_C2,
         P1_N111, P1_N110, P1_N109, P1_N108, P1_N107, P1_N106, P1_N105,
         P1_N104, P2_N111, P2_N110, P2_N109, P2_N108, P2_N107, P2_N106,
         P2_N105, P2_N104, C1_stall, C1_addr_0_, C1_addr_1_, C1_addr_2_,
         C1_addr_3_, C1_addr_4_, C1_addr_5_, C1_addr_6_, C1_addr_7_,
         C1_addr_8_, C1_addr_9_, C1_addr_10_, C1_addr_14_, C1_addr_15_, C1_N80,
         C2_stall, C2_addr_0_, C2_addr_2_, C2_addr_4_, C2_addr_5_, C2_addr_6_,
         C2_addr_7_, C2_addr_8_, C2_addr_9_, C2_addr_10_, C2_addr_11_,
         C2_addr_12_, C2_addr_13_, C2_addr_14_, C2_addr_15_, mb_stall,
         mb_prefer, mb_chipSelect, n142, n146, n147, n148, n150, n151, n155,
         n157, n159, n160, n161, n414, n416, n417, n418, n420, n424, n425,
         n431, n435, n436, n437, n438, n439, n440, n441, n442, n444, n447,
         n449, n456, n463, n464, n465, n495, n496, n500, n501, n510, n511,
         n513, n522, n527, n528, n529, n534, n536, n537, n538, n539, n542,
         n543, n547, n548, n550, n551, n552, n553, n554, n555, n556, n560,
         n561, n564, n565, n569, n570, n571, n574, n575, n577, n583, n584,
         n587, n591, n592, n600, n604, n624, n630, n631, n639, n640, n641,
         n649, n650, n652, n653, n654, n655, n656, n657, n658, n659, n662,
         n663, n664, n666, n667, n671, n672, n673, n681, n683, n685, n686,
         n689, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n707, n708, n709, n710, n711, n712, n713, n716, n719, n721,
         n722, n723, n724, n725, n729, n731, n732, n736, n737, n801, n872,
         n873, n874, n931, n932, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1228, n1250,
         n1274, n1276, n1277, n1278, n1279, n1280, n1281, n1284, n1285, n1290,
         n1293, n1294, n1296, n1297, n1359, n1404, n1405, n1407, n1408, n1409,
         n1410, n1411, n1416, n1417, n1418, n1419, n1424, n1425, n1426, n1427,
         n1432, n1433, n1434, n1438, n1441, n1442, n1444, n1445, n1446, n1448,
         n1450, n1451, n1452, n1454, n1455, n1456, n1457, n1459, n1460, n1461,
         n1464, n1466, n1471, n1473, n1474, n1475, n1476, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1488, n1517, n1518, n1521,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1542, n1543, n1544,
         n1545, n1546, n1547, n1553, n1555, n1556, n1560, n1561, n1563, n1564,
         n1568, n1569, n1570, n1571, n1575, n1576, n1577, n1579, n1580, n1585,
         n1586, n1587, n1588, n1592, n1624, n1627, n1634, n1635, n1636, n1654,
         n1655, n1656, n1657, n1658, n1659, n1662, n1663, n1664, n1669, n1671,
         n1672, n1674, n1675, n1676, n1677, n1678, n1679, n1681, n1683, n1684,
         n1685, n1686, n1687, n1688, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1707, n1708, n1713, n1714, n1715, n1737, n1738, n1740,
         n1741, n1742, n1743, n1744, n1780, n1785, n1787, n1788, n1789, n1790,
         n1791, n1792, n1801, n1802, n1804, n1811, n1812, n1817, n1818, n1819,
         n1840, n1842, n1843, n1844, n1849, n1855, n1857, n1865, n1866, n1870,
         n1871, n1898, n1901, n1916, n2011, n2389, n2391, n2394, n2395, n2403,
         n2407, n2411, n2412, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2509, n2512,
         n2514, n2515, n2516, n2521, n2522, n2523, n2524, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2538, n2539, n2540, n2541, n2542, n2545,
         n2546, n2549, n2550, n2551, n2555, n2556, n2557, n2558, n2559, n2560,
         n2562, n2563, n2564, n2570, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100;
  wire   [1:0] rw_P1_C1;
  wire   [15:0] addr_P1_C1;
  wire   [1:0] stateP1;
  wire   [1:0] rw_P2_C2;
  wire   [15:0] addr_P2_C2;
  wire   [1:0] stateP2;
  wire   [1:0] rw_C1_M;
  wire   [15:0] addr_C1_M;
  wire   [15:0] allowReadAddr_C2_C1;
  wire   [15:0] addr_C2_C1;
  wire   [15:0] allowReadAddr_C1_C2;
  wire   [15:0] addr_C1_C2;
  wire   [3:0] debugStateC1;
  wire   [1:0] rw_C2_M;
  wire   [15:0] addr_C2_M;
  wire   [3:0] debugStateC2;
  wire   [1:0] debugRwToMem;
  wire   [6:0] debugDelay;

  LVT_OAI21HSV2 U47 ( .A1(n440), .A2(n441), .B(n438), .ZN(n439) );
  LVT_INOR2HSV4 U48 ( .A1(n442), .B1(reset), .ZN(n438) );
  LVT_OAI21HSV2 U92 ( .A1(reset), .A2(n495), .B(n496), .ZN(n1074) );
  LVT_AO22HSV0 U141 ( .A1(pc_proc2_code2[6]), .A2(n550), .B1(P2_N110), .B2(
        n551), .Z(n1094) );
  LVT_AO22HSV0 U142 ( .A1(pc_proc2_code2[5]), .A2(n550), .B1(P2_N109), .B2(
        n551), .Z(n1095) );
  LVT_AO22HSV0 U143 ( .A1(pc_proc2_code2[4]), .A2(n550), .B1(P2_N108), .B2(
        n551), .Z(n1096) );
  LVT_AO22HSV0 U144 ( .A1(pc_proc2_code2[3]), .A2(n550), .B1(P2_N107), .B2(
        n551), .Z(n1097) );
  LVT_AO22HSV0 U145 ( .A1(pc_proc2_code2[2]), .A2(n550), .B1(P2_N106), .B2(
        n551), .Z(n1098) );
  LVT_AO22HSV0 U146 ( .A1(pc_proc2_code2[1]), .A2(n550), .B1(P2_N105), .B2(
        n551), .Z(n1099) );
  LVT_AO22HSV0 U147 ( .A1(pc_proc2_code2[0]), .A2(n550), .B1(P2_N104), .B2(
        n551), .Z(n1100) );
  LVT_AO22HSV0 U148 ( .A1(pc_proc2_code2[7]), .A2(n550), .B1(P2_N111), .B2(
        n551), .Z(n1101) );
  LVT_OAI32HSV2 U178 ( .A1(n574), .A2(reset), .A3(n150), .B1(n2464), .B2(n575), 
        .ZN(n1106) );
  LVT_AO22HSV0 U257 ( .A1(pc_proc1_code1[6]), .A2(n652), .B1(P1_N110), .B2(
        n653), .Z(n1144) );
  LVT_AO22HSV0 U258 ( .A1(pc_proc1_code1[5]), .A2(n652), .B1(P1_N109), .B2(
        n653), .Z(n1145) );
  LVT_AO22HSV0 U259 ( .A1(pc_proc1_code1[4]), .A2(n652), .B1(P1_N108), .B2(
        n653), .Z(n1146) );
  LVT_AO22HSV0 U260 ( .A1(pc_proc1_code1[3]), .A2(n652), .B1(P1_N107), .B2(
        n653), .Z(n1147) );
  LVT_AO22HSV0 U261 ( .A1(pc_proc1_code1[2]), .A2(n652), .B1(P1_N106), .B2(
        n653), .Z(n1148) );
  LVT_AO22HSV0 U262 ( .A1(pc_proc1_code1[1]), .A2(n652), .B1(P1_N105), .B2(
        n653), .Z(n1149) );
  LVT_AO22HSV0 U263 ( .A1(pc_proc1_code1[0]), .A2(n652), .B1(P1_N104), .B2(
        n653), .Z(n1150) );
  LVT_AO22HSV0 U264 ( .A1(pc_proc1_code1[7]), .A2(n652), .B1(P1_N111), .B2(
        n653), .Z(n1151) );
  LVT_OAI31HSV2 U273 ( .A1(n666), .A2(n662), .A3(n2589), .B(n658), .ZN(n664)
         );
  LVT_OAI222HSV2 U310 ( .A1(n3091), .A2(n695), .B1(n2532), .B2(n696), .C1(n697), .C2(n2450), .ZN(n1160) );
  LVT_OAI222HSV2 U312 ( .A1(n3093), .A2(n695), .B1(n2516), .B2(n696), .C1(n697), .C2(n2441), .ZN(n1162) );
  LVT_OAI222HSV2 U313 ( .A1(n3094), .A2(n695), .B1(n2515), .B2(n696), .C1(n697), .C2(n2447), .ZN(n1163) );
  LVT_OAI222HSV2 U317 ( .A1(n3087), .A2(n695), .B1(n2523), .B2(n696), .C1(n697), .C2(n2448), .ZN(n1167) );
  LVT_OAI222HSV2 U320 ( .A1(n3095), .A2(n695), .B1(n2564), .B2(n696), .C1(n697), .C2(n2427), .ZN(n1170) );
  LVT_OAI222HSV2 U321 ( .A1(n3089), .A2(n695), .B1(n1285), .B2(n696), .C1(n697), .C2(n2416), .ZN(n1171) );
  LVT_OAI21HSV2 U349 ( .A1(n721), .A2(n722), .B(n723), .ZN(n1187) );
  LVT_OAI21HSV2 U350 ( .A1(n3047), .A2(n721), .B(allowRead_C2_C1), .ZN(n723)
         );
  LVT_OAI222HSV2 U453 ( .A1(n3085), .A2(n695), .B1(n2534), .B2(n696), .C1(n697), .C2(n2439), .ZN(n1191) );
  LVT_OAI21HSV2 U458 ( .A1(n3037), .A2(n732), .B(n801), .ZN(n695) );
  LVT_OAI222HSV2 U567 ( .A1(n2509), .A2(n872), .B1(n2545), .B2(n873), .C1(n874), .C2(n2475), .ZN(n1192) );
  LVT_OAI222HSV2 U568 ( .A1(n2575), .A2(n872), .B1(n1281), .B2(n873), .C1(n874), .C2(n2476), .ZN(n1193) );
  LVT_OAI222HSV2 U569 ( .A1(n2574), .A2(n872), .B1(n1297), .B2(n873), .C1(n874), .C2(n2487), .ZN(n1194) );
  LVT_OAI222HSV2 U570 ( .A1(n2576), .A2(n872), .B1(n1279), .B2(n873), .C1(n874), .C2(n2473), .ZN(n1195) );
  LVT_OAI222HSV2 U571 ( .A1(n2529), .A2(n872), .B1(n2524), .B2(n873), .C1(n874), .C2(n2490), .ZN(n1196) );
  LVT_OAI222HSV2 U572 ( .A1(n2531), .A2(n872), .B1(n2521), .B2(n873), .C1(n874), .C2(n2491), .ZN(n1197) );
  LVT_OAI222HSV2 U573 ( .A1(n2530), .A2(n872), .B1(n2541), .B2(n873), .C1(n874), .C2(n2470), .ZN(n1198) );
  LVT_OAI222HSV2 U574 ( .A1(n2514), .A2(n872), .B1(n2522), .B2(n873), .C1(n874), .C2(n2471), .ZN(n1199) );
  LVT_OAI222HSV2 U575 ( .A1(n2557), .A2(n872), .B1(n2538), .B2(n873), .C1(n874), .C2(n2481), .ZN(n1200) );
  LVT_OAI222HSV2 U576 ( .A1(n2550), .A2(n872), .B1(n2542), .B2(n873), .C1(n874), .C2(n2496), .ZN(n1201) );
  LVT_OAI222HSV2 U577 ( .A1(n2578), .A2(n872), .B1(n2579), .B2(n873), .C1(n874), .C2(n2480), .ZN(n1202) );
  LVT_OAI222HSV2 U578 ( .A1(n2581), .A2(n872), .B1(n2540), .B2(n873), .C1(n874), .C2(n2502), .ZN(n1203) );
  LVT_OAI222HSV2 U579 ( .A1(n2549), .A2(n872), .B1(n2539), .B2(n873), .C1(n874), .C2(n2506), .ZN(n1204) );
  LVT_OAI222HSV2 U580 ( .A1(n2551), .A2(n872), .B1(n2555), .B2(n873), .C1(n874), .C2(n2507), .ZN(n1205) );
  LVT_OAI222HSV2 U593 ( .A1(n2577), .A2(n872), .B1(n2580), .B2(n873), .C1(n874), .C2(n2486), .ZN(n1208) );
  LVT_OAI21HSV2 U714 ( .A1(n3064), .A2(n600), .B(C1_N80), .ZN(n604) );
  LVT_OAI32HSV2 U791 ( .A1(n159), .A2(mb_chipSelect), .A3(n155), .B1(n3064), 
        .B2(n698), .ZN(n1210) );
  LVT_OAI21HSV2 U800 ( .A1(n711), .A2(n712), .B(n1870), .ZN(n1018) );
  LVT_CLKNHSV2 U805 ( .I(reset), .ZN(C1_N80) );
  LVT_CLKNHSV2 U807 ( .I(n584), .ZN(n142) );
  LVT_CLKNHSV2 U811 ( .I(n686), .ZN(n146) );
  LVT_CLKNHSV2 U822 ( .I(n1018), .ZN(n157) );
  LVT_CLKNHSV2 U824 ( .I(n699), .ZN(n159) );
  LVT_CLKNHSV2 U825 ( .I(n658), .ZN(n160) );
  LVT_CLKNHSV2 U826 ( .I(n556), .ZN(n161) );
  LVT_DQHSV1 C2_addrToCache_reg_14_ ( .D(n1038), .CK(clk), .Q(addr_C2_C1[14])
         );
  LVT_DQHSV1 C2_addrToCache_reg_13_ ( .D(n1039), .CK(clk), .Q(addr_C2_C1[13])
         );
  LVT_DQHSV1 C1_addrToMem_reg_0_ ( .D(n1122), .CK(clk), .Q(addr_C1_M[0]) );
  LVT_DQHSV1 C2_addrToMem_reg_1_ ( .D(n1171), .CK(clk), .Q(addr_C2_M[1]) );
  LVT_DQHSV1 C1_addrToMem_reg_14_ ( .D(n1108), .CK(clk), .Q(addr_C1_M[14]) );
  LVT_DQHSV1 C1_addrToMem_reg_13_ ( .D(n1109), .CK(clk), .Q(addr_C1_M[13]) );
  LVT_DQHSV1 C1_addrToMem_reg_12_ ( .D(n1110), .CK(clk), .Q(addr_C1_M[12]) );
  LVT_DQHSV1 C1_addrToMem_reg_8_ ( .D(n1114), .CK(clk), .Q(addr_C1_M[8]) );
  LVT_DQHSV1 C1_addrToMem_reg_4_ ( .D(n1118), .CK(clk), .Q(addr_C1_M[4]) );
  LVT_DQHSV1 C1_addrToMem_reg_3_ ( .D(n1119), .CK(clk), .Q(addr_C1_M[3]) );
  LVT_DQHSV1 C1_addrToMem_reg_2_ ( .D(n1120), .CK(clk), .Q(addr_C1_M[2]) );
  LVT_DQHSV1 C1_addrToMem_reg_1_ ( .D(n1121), .CK(clk), .Q(addr_C1_M[1]) );
  LVT_DQHSV1 C1_addrToMem_reg_15_ ( .D(n1207), .CK(clk), .Q(addr_C1_M[15]) );
  LVT_DQHSV1 C2_addrToMem_reg_3_ ( .D(n1169), .CK(clk), .Q(addr_C2_M[3]) );
  LVT_DQHSV1 C2_addrToMem_reg_2_ ( .D(n1170), .CK(clk), .Q(addr_C2_M[2]) );
  LVT_DQHSV1 C1_addrToMem_reg_11_ ( .D(n1111), .CK(clk), .Q(addr_C1_M[11]) );
  LVT_DQHSV1 C1_addrToMem_reg_10_ ( .D(n1112), .CK(clk), .Q(addr_C1_M[10]) );
  LVT_DQHSV1 C1_addrToMem_reg_9_ ( .D(n1113), .CK(clk), .Q(addr_C1_M[9]) );
  LVT_DQHSV1 C1_addrToMem_reg_7_ ( .D(n1115), .CK(clk), .Q(addr_C1_M[7]) );
  LVT_DQHSV1 C1_addrToMem_reg_6_ ( .D(n1116), .CK(clk), .Q(addr_C1_M[6]) );
  LVT_DQHSV1 C1_addrToMem_reg_5_ ( .D(n1117), .CK(clk), .Q(addr_C1_M[5]) );
  LVT_DQHSV1 mb_delay_reg_4_ ( .D(n1179), .CK(clk), .Q(debugDelay[4]) );
  LVT_DQHSV1 C1_addrToCache_reg_7_ ( .D(n1064), .CK(clk), .Q(addr_C1_C2[7]) );
  LVT_DQHSV1 C1_addrToCache_reg_14_ ( .D(n1057), .CK(clk), .Q(addr_C1_C2[14])
         );
  LVT_DQHSV1 C1_addrToCache_reg_10_ ( .D(n1061), .CK(clk), .Q(addr_C1_C2[10])
         );
  LVT_DQHSV1 C1_addrToCache_reg_6_ ( .D(n1065), .CK(clk), .Q(addr_C1_C2[6]) );
  LVT_DQHSV1 C1_addrToCache_reg_11_ ( .D(n1060), .CK(clk), .Q(addr_C1_C2[11])
         );
  LVT_DQHSV1 C1_addrToCache_reg_4_ ( .D(n1067), .CK(clk), .Q(addr_C1_C2[4]) );
  LVT_DQHSV1 C1_addrToCache_reg_5_ ( .D(n1066), .CK(clk), .Q(addr_C1_C2[5]) );
  LVT_DQHSV1 C1_rwToMem_reg_1_ ( .D(n1186), .CK(clk), .Q(rw_C1_M[1]) );
  LVT_DQHSV1 C1_wmToCache_reg ( .D(n1072), .CK(clk), .Q(wm_C1_C2) );
  LVT_DQHSV1 C2_addrToMem_reg_0_ ( .D(n1172), .CK(clk), .Q(addr_C2_M[0]) );
  LVT_DQHSV1 C2_addrToCache_reg_0_ ( .D(n1052), .CK(clk), .Q(addr_C2_C1[0]) );
  LVT_DQHSV1 C2_addrToMem_reg_15_ ( .D(n1191), .CK(clk), .Q(addr_C2_M[15]) );
  LVT_DQHSV1 C2_addrToMem_reg_8_ ( .D(n1164), .CK(clk), .Q(addr_C2_M[8]) );
  LVT_DQHSV1 C2_addrToMem_reg_10_ ( .D(n1162), .CK(clk), .Q(addr_C2_M[10]) );
  LVT_DQHSV1 C2_addrToMem_reg_7_ ( .D(n1165), .CK(clk), .Q(addr_C2_M[7]) );
  LVT_DQHSV1 C2_addrToMem_reg_6_ ( .D(n1166), .CK(clk), .Q(addr_C2_M[6]) );
  LVT_DQHSV1 C2_addrToMem_reg_4_ ( .D(n1168), .CK(clk), .Q(addr_C2_M[4]) );
  LVT_DQHSV1 C2_addrToMem_reg_13_ ( .D(n1159), .CK(clk), .Q(addr_C2_M[13]) );
  LVT_DQHSV1 C2_addrToMem_reg_11_ ( .D(n1161), .CK(clk), .Q(addr_C2_M[11]) );
  LVT_DQHSV1 C2_addrToMem_reg_9_ ( .D(n1163), .CK(clk), .Q(addr_C2_M[9]) );
  LVT_DQHSV1 C2_addrToMem_reg_5_ ( .D(n1167), .CK(clk), .Q(addr_C2_M[5]) );
  LVT_DQHSV1 C2_addrToMem_reg_14_ ( .D(n1158), .CK(clk), .Q(addr_C2_M[14]) );
  LVT_DQHSV1 C2_addrToMem_reg_12_ ( .D(n1160), .CK(clk), .Q(addr_C2_M[12]) );
  LVT_DQHSV1 mb_delay_reg_2_ ( .D(n1181), .CK(clk), .Q(debugDelay[2]) );
  LVT_DQHSV1 C1_addrToCache_reg_1_ ( .D(n1070), .CK(clk), .Q(addr_C1_C2[1]) );
  LVT_DQHSV1 mb_delay_reg_1_ ( .D(n1182), .CK(clk), .Q(debugDelay[1]) );
  LVT_DQHSV1 C2_rmToCache_reg ( .D(n1157), .CK(clk), .Q(rm_C2_C1) );
  LVT_DQHSV1 C1_addrToCache_reg_15_ ( .D(n1056), .CK(clk), .Q(addr_C1_C2[15])
         );
  LVT_DQHSV1 C1_havMsgToCache_reg ( .D(n1055), .CK(clk), .Q(msg_C1_C2) );
  LVT_DQHSV1 mb_prefer_reg ( .D(n1175), .CK(clk), .Q(mb_prefer) );
  LVT_DQHSV1 P1_rwToMem_reg_1_ ( .D(n1152), .CK(clk), .Q(rw_P1_C1[1]) );
  LVT_DQHSV1 C2_rwToMem_reg_0_ ( .D(n1019), .CK(clk), .Q(rw_C2_M[0]) );
  LVT_DQHSV1 C1_addrToCache_reg_0_ ( .D(n1071), .CK(clk), .Q(addr_C1_C2[0]) );
  LVT_DQHSV1 C1_addrToCache_reg_2_ ( .D(n1069), .CK(clk), .Q(addr_C1_C2[2]) );
  LVT_DQHSV1 C1_allowReadToCache_reg ( .D(n1188), .CK(clk), .Q(allowRead_C1_C2) );
  LVT_DQHSV1 mb_rwToMem_reg_0_ ( .D(n1184), .CK(clk), .Q(debugRwToMem[0]) );
  LVT_DQHSV1 C1_rwToMem_reg_0_ ( .D(n1123), .CK(clk), .Q(rw_C1_M[0]) );
  LVT_DQHSV1 C2_addrToCache_reg_4_ ( .D(n1048), .CK(clk), .Q(addr_C2_C1[4]) );
  LVT_DQHSV1 C2_addrToCache_reg_8_ ( .D(n1044), .CK(clk), .Q(addr_C2_C1[8]) );
  LVT_DQHSV1 C2_addrToCache_reg_15_ ( .D(n1037), .CK(clk), .Q(addr_C2_C1[15])
         );
  LVT_DQHSV1 C2_addrToCache_reg_3_ ( .D(n1049), .CK(clk), .Q(addr_C2_C1[3]) );
  LVT_DQHSV1 C2_addrToCache_reg_2_ ( .D(n1050), .CK(clk), .Q(addr_C2_C1[2]) );
  LVT_DQHSV1 C2_addrToCache_reg_1_ ( .D(n1051), .CK(clk), .Q(addr_C2_C1[1]) );
  LVT_DQHSV1 mb_chipSelect_reg ( .D(n1211), .CK(clk), .Q(mb_chipSelect) );
  LVT_DQHSV1 C2_cacheEnToCPU_reg ( .D(n1106), .CK(clk), .Q(en_C2_P2) );
  LVT_DQHSV1 C1_cacheEnToCPU_reg ( .D(n1156), .CK(clk), .Q(en_C1_P1) );
  LVT_DQHSV1 mb_delay_reg_0_ ( .D(n1183), .CK(clk), .Q(debugDelay[0]) );
  LVT_DQHSV1 P2_state_reg_1_ ( .D(n1105), .CK(clk), .Q(stateP2[1]) );
  LVT_DQHSV1 C2_stall_reg ( .D(n1021), .CK(clk), .Q(C2_stall) );
  LVT_DQHSV1 P1_state_reg_1_ ( .D(n1155), .CK(clk), .Q(stateP1[1]) );
  LVT_DQHSV1 C2_addrToCache_reg_5_ ( .D(n1047), .CK(clk), .Q(addr_C2_C1[5]) );
  LVT_DQHSV1 C2_addrToCache_reg_9_ ( .D(n1043), .CK(clk), .Q(addr_C2_C1[9]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_8_ ( .D(n1028), .CK(clk), .Q(
        allowReadAddr_C2_C1[8]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_7_ ( .D(n1029), .CK(clk), .Q(
        allowReadAddr_C2_C1[7]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_8_ ( .D(n1198), .CK(clk), .Q(
        allowReadAddr_C1_C2[8]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_7_ ( .D(n1199), .CK(clk), .Q(
        allowReadAddr_C1_C2[7]) );
  LVT_DQHSV1 C2_havMsgToCache_reg ( .D(n1074), .CK(clk), .Q(msg_C2_C1) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_11_ ( .D(n1025), .CK(clk), .Q(
        allowReadAddr_C2_C1[11]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_11_ ( .D(n1195), .CK(clk), .Q(
        allowReadAddr_C1_C2[11]) );
  LVT_DQHSV1 mb_stall_reg ( .D(n1174), .CK(clk), .Q(mb_stall) );
  LVT_DQHSV1 C2_allowReadToCache_reg ( .D(n1187), .CK(clk), .Q(allowRead_C2_C1) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_14_ ( .D(n1192), .CK(clk), .Q(
        allowReadAddr_C1_C2[14]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_13_ ( .D(n1193), .CK(clk), .Q(
        allowReadAddr_C1_C2[13]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_3_ ( .D(n1033), .CK(clk), .Q(
        allowReadAddr_C2_C1[3]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_4_ ( .D(n1032), .CK(clk), .Q(
        allowReadAddr_C2_C1[4]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_6_ ( .D(n1030), .CK(clk), .Q(
        allowReadAddr_C2_C1[6]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_4_ ( .D(n1202), .CK(clk), .Q(
        allowReadAddr_C1_C2[4]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_6_ ( .D(n1200), .CK(clk), .Q(
        allowReadAddr_C1_C2[6]) );
  LVT_DQHSV1 C1_rmToCache_reg ( .D(n1107), .CK(clk), .Q(rm_C1_C2) );
  LVT_DQHSV1 C1_stall_reg ( .D(n1124), .CK(clk), .Q(C1_stall) );
  LVT_DQHSV1 C2_wmToCache_reg ( .D(n1053), .CK(clk), .Q(wm_C2_C1) );
  LVT_DQHSV1 mb_delay_reg_6_ ( .D(n1177), .CK(clk), .Q(debugDelay[6]) );
  LVT_DQHSV1 mb_delay_reg_3_ ( .D(n1180), .CK(clk), .Q(debugDelay[3]) );
  LVT_DQHSV1 C2_rwToMem_reg_1_ ( .D(n1020), .CK(clk), .Q(rw_C2_M[1]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_15_ ( .D(n1208), .CK(clk), .Q(
        allowReadAddr_C1_C2[15]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_12_ ( .D(n1194), .CK(clk), .Q(
        allowReadAddr_C1_C2[12]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_10_ ( .D(n1026), .CK(clk), .Q(
        allowReadAddr_C2_C1[10]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_9_ ( .D(n1027), .CK(clk), .Q(
        allowReadAddr_C2_C1[9]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_10_ ( .D(n1196), .CK(clk), .Q(
        allowReadAddr_C1_C2[10]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_9_ ( .D(n1197), .CK(clk), .Q(
        allowReadAddr_C1_C2[9]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_2_ ( .D(n1034), .CK(clk), .Q(
        allowReadAddr_C2_C1[2]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_1_ ( .D(n1035), .CK(clk), .Q(
        allowReadAddr_C2_C1[1]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_5_ ( .D(n1031), .CK(clk), .Q(
        allowReadAddr_C2_C1[5]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_0_ ( .D(n1036), .CK(clk), .Q(
        allowReadAddr_C2_C1[0]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_5_ ( .D(n1201), .CK(clk), .Q(
        allowReadAddr_C1_C2[5]) );
  LVT_DQHSV1 P2_addrToMem_reg_1_ ( .D(n1092), .CK(clk), .Q(addr_P2_C2[1]) );
  LVT_DQHSV1 P1_state_reg_0_ ( .D(n1154), .CK(clk), .Q(stateP1[0]) );
  LVT_DQHSV1 mb_rwToMem_reg_1_ ( .D(n1185), .CK(clk), .Q(debugRwToMem[1]) );
  LVT_DQHSV1 P2_addrToMem_reg_2_ ( .D(n1091), .CK(clk), .Q(addr_P2_C2[2]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_12_ ( .D(n1024), .CK(clk), .Q(
        allowReadAddr_C2_C1[12]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_0_ ( .D(n1206), .CK(clk), .Q(
        allowReadAddr_C1_C2[0]) );
  LVT_DQHSV1 mb_delay_reg_5_ ( .D(n1178), .CK(clk), .Q(debugDelay[5]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_3_ ( .D(n1203), .CK(clk), .Q(
        allowReadAddr_C1_C2[3]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_15_ ( .D(n1189), .CK(clk), .Q(
        allowReadAddr_C2_C1[15]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_14_ ( .D(n1022), .CK(clk), .Q(
        allowReadAddr_C2_C1[14]) );
  LVT_DQHSV1 C2_allowReadToCacheAddr_reg_13_ ( .D(n1023), .CK(clk), .Q(
        allowReadAddr_C2_C1[13]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_2_ ( .D(n1204), .CK(clk), .Q(
        allowReadAddr_C1_C2[2]) );
  LVT_DQHSV1 C1_allowReadToCacheAddr_reg_1_ ( .D(n1205), .CK(clk), .Q(
        allowReadAddr_C1_C2[1]) );
  LVT_DQHSV1 P2_state_reg_0_ ( .D(n1104), .CK(clk), .Q(stateP2[0]) );
  LVT_DQHSV1 P1_addrToMem_reg_14_ ( .D(n1129), .CK(clk), .Q(addr_P1_C1[14]) );
  LVT_DQHSV1 P1_counter_reg_7_ ( .D(n1151), .CK(clk), .Q(pc_proc1_code1[7]) );
  LVT_DQHSV1 P2_counter_reg_7_ ( .D(n1101), .CK(clk), .Q(pc_proc2_code2[7]) );
  LVT_DQHSV1 P1_rwToMem_reg_0_ ( .D(n1153), .CK(clk), .Q(rw_P1_C1[0]) );
  LVT_DQHSV1 P1_counter_reg_1_ ( .D(n1149), .CK(clk), .Q(pc_proc1_code1[1]) );
  LVT_DQHSV1 P1_counter_reg_2_ ( .D(n1148), .CK(clk), .Q(pc_proc1_code1[2]) );
  LVT_DQHSV1 P1_counter_reg_3_ ( .D(n1147), .CK(clk), .Q(pc_proc1_code1[3]) );
  LVT_DQHSV1 P1_counter_reg_4_ ( .D(n1146), .CK(clk), .Q(pc_proc1_code1[4]) );
  LVT_DQHSV1 P1_counter_reg_5_ ( .D(n1145), .CK(clk), .Q(pc_proc1_code1[5]) );
  LVT_DQHSV1 P1_counter_reg_6_ ( .D(n1144), .CK(clk), .Q(pc_proc1_code1[6]) );
  LVT_DQHSV1 P2_counter_reg_1_ ( .D(n1099), .CK(clk), .Q(pc_proc2_code2[1]) );
  LVT_DQHSV1 P2_counter_reg_2_ ( .D(n1098), .CK(clk), .Q(pc_proc2_code2[2]) );
  LVT_DQHSV1 P2_counter_reg_3_ ( .D(n1097), .CK(clk), .Q(pc_proc2_code2[3]) );
  LVT_DQHSV1 P2_counter_reg_4_ ( .D(n1096), .CK(clk), .Q(pc_proc2_code2[4]) );
  LVT_DQHSV1 P2_counter_reg_5_ ( .D(n1095), .CK(clk), .Q(pc_proc2_code2[5]) );
  LVT_DQHSV1 P2_counter_reg_6_ ( .D(n1094), .CK(clk), .Q(pc_proc2_code2[6]) );
  LVT_DQHSV1 P1_counter_reg_0_ ( .D(n1150), .CK(clk), .Q(pc_proc1_code1[0]) );
  LVT_DQHSV1 P2_counter_reg_0_ ( .D(n1100), .CK(clk), .Q(pc_proc2_code2[0]) );
  LVT_DQHSV1 P2_addrToMem_reg_5_ ( .D(n1088), .CK(clk), .Q(addr_P2_C2[5]) );
  LVT_DQHSV1 P1_addrToMem_reg_7_ ( .D(n1136), .CK(clk), .Q(addr_P1_C1[7]) );
  LVT_DQHSV1 P2_rwToMem_reg_0_ ( .D(n1103), .CK(clk), .Q(rw_P2_C2[0]) );
  HVT_DQHSV1 P2_rwToMem_reg_1_ ( .D(n1102), .CK(clk), .Q(rw_P2_C2[1]) );
  LVT_EDGRNQHSV1 C1_addr_reg_7_ ( .RN(C1_N80), .D(addr_C1_M[7]), .E(n2951), 
        .CK(clk), .Q(C1_addr_7_) );
  LVT_DQHSV1 P2_addrToMem_reg_15_ ( .D(n1078), .CK(clk), .Q(addr_P2_C2[15]) );
  LVT_DQHSV1 P2_addrToMem_reg_11_ ( .D(n1082), .CK(clk), .Q(addr_P2_C2[11]) );
  LVT_DQHSV1 P2_addrToMem_reg_9_ ( .D(n1084), .CK(clk), .Q(addr_P2_C2[9]) );
  LVT_DQHSV1 P1_addrToMem_reg_10_ ( .D(n1133), .CK(clk), .Q(addr_P1_C1[10]) );
  LVT_DQHSV1 P1_addrToMem_reg_8_ ( .D(n1135), .CK(clk), .Q(addr_P1_C1[8]) );
  LVT_DQHSV1 P1_addrToMem_reg_9_ ( .D(n1134), .CK(clk), .Q(addr_P1_C1[9]) );
  LVT_EDGRNQHSV1 C1_addr_reg_6_ ( .RN(C1_N80), .D(addr_C1_M[6]), .E(n3031), 
        .CK(clk), .Q(C1_addr_6_) );
  LVT_EDGRNQHSV1 C1_addr_reg_2_ ( .RN(C1_N80), .D(addr_C1_M[2]), .E(n2951), 
        .CK(clk), .Q(C1_addr_2_) );
  LVT_EDGRNQHSV1 C1_addr_reg_3_ ( .RN(C1_N80), .D(addr_C1_M[3]), .E(n3030), 
        .CK(clk), .Q(C1_addr_3_) );
  LVT_EDGRNQHSV1 C1_addr_reg_8_ ( .RN(C1_N80), .D(addr_C1_M[8]), .E(n2951), 
        .CK(clk), .Q(C1_addr_8_) );
  LVT_EDGRNQHSV1 C1_addr_reg_5_ ( .RN(C1_N80), .D(addr_C1_M[5]), .E(n3030), 
        .CK(clk), .Q(C1_addr_5_) );
  LVT_EDGRNQHSV1 C1_addr_reg_0_ ( .RN(C1_N80), .D(addr_C1_M[0]), .E(n3031), 
        .CK(clk), .Q(C1_addr_0_) );
  LVT_EDGRNQHSV1 C1_addr_reg_14_ ( .RN(C1_N80), .D(addr_C1_M[14]), .E(n3030), 
        .CK(clk), .Q(C1_addr_14_) );
  LVT_DQHSV1 C1_addrToCache_reg_12_ ( .D(n1059), .CK(clk), .Q(addr_C1_C2[12])
         );
  LVT_DQHSV1 C1_addrToCache_reg_13_ ( .D(n1058), .CK(clk), .Q(addr_C1_C2[13])
         );
  LVT_DQHSV1 P1_addrToMem_reg_2_ ( .D(n1141), .CK(clk), .Q(addr_P1_C1[2]) );
  LVT_DQHSV1 P1_addrToMem_reg_5_ ( .D(n1138), .CK(clk), .Q(addr_P1_C1[5]) );
  LVT_DQHSV1 P1_addrToMem_reg_1_ ( .D(n1142), .CK(clk), .Q(addr_P1_C1[1]) );
  LVT_DQHSV1 P1_addrToMem_reg_0_ ( .D(n1143), .CK(clk), .Q(addr_P1_C1[0]) );
  LVT_DQHSV1 C1_addrToCache_reg_9_ ( .D(n1062), .CK(clk), .Q(addr_C1_C2[9]) );
  LVT_DQHSV1 C1_addrToCache_reg_3_ ( .D(n1068), .CK(clk), .Q(addr_C1_C2[3]) );
  LVT_DQHSV1 C1_addrToCache_reg_8_ ( .D(n1063), .CK(clk), .Q(addr_C1_C2[8]) );
  LVT_EDGRNQHSV1 C1_addr_reg_1_ ( .RN(C1_N80), .D(addr_C1_M[1]), .E(n3031), 
        .CK(clk), .Q(C1_addr_1_) );
  LVT_DQHSV1 C2_addrToCache_reg_11_ ( .D(n1041), .CK(clk), .Q(addr_C2_C1[11])
         );
  LVT_DQHSV1 P1_addrToMem_reg_6_ ( .D(n1137), .CK(clk), .Q(addr_P1_C1[6]) );
  LVT_DQHSV1 C2_addrToCache_reg_7_ ( .D(n1045), .CK(clk), .Q(addr_C2_C1[7]) );
  LVT_DQHSV1 C2_addrToCache_reg_6_ ( .D(n1046), .CK(clk), .Q(addr_C2_C1[6]) );
  LVT_EDGRNHSV1 C1_addr_reg_12_ ( .RN(C1_N80), .D(addr_C1_M[12]), .E(n3031), 
        .CK(clk), .Q(n1296), .QN(n1297) );
  LVT_DHSV1 C2_addrToCache_reg_10_ ( .D(n1042), .CK(clk), .Q(n1293), .QN(n1294) );
  LVT_DQHSV1 C2_addrToCache_reg_12_ ( .D(n1040), .CK(clk), .Q(addr_C2_C1[12])
         );
  LVT_DQHSV1 P2_addrToMem_reg_6_ ( .D(n1087), .CK(clk), .Q(addr_P2_C2[6]) );
  HVT_AO22HSV1 U1067 ( .A1(n1659), .A2(addr_P1_C1[2]), .B1(addr_C1_C2[2]), 
        .B2(n1658), .Z(n1069) );
  HVT_AO22HSV1 U1080 ( .A1(n1659), .A2(addr_P1_C1[11]), .B1(addr_C1_C2[11]), 
        .B2(n1658), .Z(n1060) );
  HVT_AO22HSV1 U1082 ( .A1(n1659), .A2(addr_P1_C1[13]), .B1(addr_C1_C2[13]), 
        .B2(n1658), .Z(n1058) );
  HVT_AO22HSV1 U1084 ( .A1(n1659), .A2(addr_P1_C1[12]), .B1(addr_C1_C2[12]), 
        .B2(n1658), .Z(n1059) );
  LVT_OAI211HSV4 U1104 ( .A1(n3049), .A2(n1635), .B(n1818), .C(n1707), .ZN(
        n872) );
  LVT_NAND2HSV2 U1164 ( .A1(n1787), .A2(n1788), .ZN(n1359) );
  LVT_INOR2HSV4 U1169 ( .A1(n425), .B1(reset), .ZN(n801) );
  LVT_OR4HSV2 U1181 ( .A1(n3045), .A2(n1707), .A3(n604), .A4(n3036), .Z(n1708)
         );
  LVT_AND2HSV4 U1192 ( .A1(n725), .A2(C1_N80), .Z(n731) );
  LVT_OAI221HSV1 U1246 ( .A1(n537), .A2(n534), .B1(en_M_C2), .B2(n538), .C(
        n539), .ZN(n527) );
  LVT_OAI222HSV0 U1249 ( .A1(n3085), .A2(n435), .B1(n2534), .B2(n436), .C1(
        n437), .C2(n2503), .ZN(n1189) );
  LVT_OAI222HSV0 U1250 ( .A1(n3091), .A2(n435), .B1(n2532), .B2(n436), .C1(
        n437), .C2(n2499), .ZN(n1024) );
  LVT_OAI222HSV0 U1251 ( .A1(n3087), .A2(n435), .B1(n2523), .B2(n436), .C1(
        n437), .C2(n2494), .ZN(n1031) );
  LVT_OAI222HSV0 U1252 ( .A1(n3089), .A2(n435), .B1(n1285), .B2(n436), .C1(
        n437), .C2(n2493), .ZN(n1035) );
  LVT_OAI222HSV0 U1253 ( .A1(n3095), .A2(n435), .B1(n2564), .B2(n436), .C1(
        n437), .C2(n2492), .ZN(n1034) );
  LVT_OAI222HSV0 U1254 ( .A1(n3094), .A2(n435), .B1(n2515), .B2(n436), .C1(
        n437), .C2(n2489), .ZN(n1027) );
  LVT_OAI222HSV0 U1255 ( .A1(n3093), .A2(n435), .B1(n2516), .B2(n436), .C1(
        n437), .C2(n2488), .ZN(n1026) );
  LVT_OAI211HSV1 U1257 ( .A1(n681), .A2(n1789), .B(n1788), .C(n1818), .ZN(
        n1790) );
  HVT_OAI222HSV0 U1264 ( .A1(n3092), .A2(n435), .B1(n3082), .B2(n436), .C1(
        n437), .C2(n2495), .ZN(n1036) );
  LVT_OAI21HSV1 U1268 ( .A1(n1840), .A2(n1274), .B(n1587), .ZN(n1019) );
  LVT_OAI222HSV0 U1362 ( .A1(n3088), .A2(n435), .B1(n3080), .B2(n436), .C1(
        n437), .C2(n2468), .ZN(n1028) );
  HVT_CLKNHSV0 U1378 ( .I(n456), .ZN(n148) );
  HVT_AO22HSV2 U1401 ( .A1(n1659), .A2(addr_P1_C1[6]), .B1(addr_C1_C2[6]), 
        .B2(n1658), .Z(n1065) );
  LVT_OAI221HSV0 U1421 ( .A1(n444), .A2(n692), .B1(n693), .B2(n694), .C(C1_N80), .ZN(n456) );
  LVT_AO22HSV1 U1423 ( .A1(n1659), .A2(addr_P1_C1[3]), .B1(addr_C1_C2[3]), 
        .B2(n1658), .Z(n1068) );
  LVT_AO22HSV1 U1424 ( .A1(n1659), .A2(addr_P1_C1[9]), .B1(addr_C1_C2[9]), 
        .B2(n1658), .Z(n1062) );
  HVT_AO22HSV0 U1426 ( .A1(addr_P1_C1[0]), .A2(n1659), .B1(addr_C1_C2[0]), 
        .B2(n1658), .Z(n1071) );
  LVT_AO22HSV1 U1427 ( .A1(n1659), .A2(addr_P1_C1[1]), .B1(addr_C1_C2[1]), 
        .B2(n1658), .Z(n1070) );
  HVT_AO22HSV1 U1429 ( .A1(n1659), .A2(addr_P1_C1[5]), .B1(addr_C1_C2[5]), 
        .B2(n1658), .Z(n1066) );
  HVT_AO22HSV1 U1430 ( .A1(n1659), .A2(addr_P1_C1[4]), .B1(addr_C1_C2[4]), 
        .B2(n1658), .Z(n1067) );
  HVT_AO22HSV2 U1437 ( .A1(n1659), .A2(addr_P1_C1[15]), .B1(addr_C1_C2[15]), 
        .B2(n1658), .Z(n1056) );
  HVT_OR3HSV2 U1462 ( .A1(n151), .A2(n1569), .A3(n3031), .Z(n1570) );
  HVT_OR3HSV1 U1463 ( .A1(n604), .A2(n3030), .A3(n3040), .Z(n1785) );
  HVT_OR3HSV1 U1464 ( .A1(n424), .A2(n3028), .A3(n425), .Z(n1585) );
  LVT_NOR4HSV0 U1476 ( .A1(n725), .A2(n577), .A3(n3046), .A4(n3071), .ZN(n721)
         );
  LVT_NAND2HSV0 U1477 ( .A1(n731), .A2(n732), .ZN(n435) );
  LVT_IOA22HSV0 U1480 ( .B1(n1857), .B2(n416), .A1(n1857), .A2(rw_C2_M[1]), 
        .ZN(n1020) );
  HVT_OAI21HSV0 U1481 ( .A1(n1555), .A2(n1801), .B(n640), .ZN(n1556) );
  LVT_INOR4HSV2 U1482 ( .A1(n587), .B1(n3036), .B2(n3042), .B3(n3060), .ZN(
        n584) );
  LVT_INOR2HSV1 U1487 ( .A1(n731), .B1(n3047), .ZN(n437) );
  LVT_NAND2HSV0 U1488 ( .A1(n731), .A2(n3035), .ZN(n436) );
  LVT_NAND2HSV0 U1498 ( .A1(n801), .A2(n3035), .ZN(n696) );
  LVT_NAND3HSV1 U1500 ( .A1(n510), .A2(n511), .A3(n3033), .ZN(n1075) );
  HVT_MUX2NHSV0 U1505 ( .I0(n1695), .I1(n3076), .S(n1697), .ZN(n1103) );
  HVT_AOI211HSV0 U1506 ( .A1(n3038), .A2(n3053), .B(n1792), .C(n1791), .ZN(
        n630) );
  LVT_NAND2HSV1 U1509 ( .A1(n931), .A2(n932), .ZN(n1209) );
  HVT_AOI211HSV0 U1510 ( .A1(n624), .A2(n465), .B(n151), .C(n464), .ZN(n931)
         );
  LVT_INOR4HSV2 U1514 ( .A1(n689), .B1(n3071), .B2(n3073), .B3(n3084), .ZN(
        n686) );
  LVT_AO32HSV0 U1515 ( .A1(n685), .A2(C1_N80), .A3(n146), .B1(n686), .B2(
        rm_C2_C1), .Z(n1157) );
  LVT_INHSV2 U1524 ( .I(n447), .ZN(n147) );
  HVT_AOI211HSV0 U1529 ( .A1(n3034), .A2(n3070), .B(n724), .C(n1901), .ZN(n722) );
  HVT_MUX2NHSV0 U1531 ( .I0(n1698), .I1(n3100), .S(n1697), .ZN(n1102) );
  LVT_AO32HSV0 U1532 ( .A1(n142), .A2(C1_N80), .A3(n583), .B1(n584), .B2(
        rm_C1_C2), .Z(n1107) );
  HVT_AOI211HSV0 U1545 ( .A1(n3038), .A2(n3043), .B(n1561), .C(n1560), .ZN(
        n1563) );
  LVT_MUX2NHSV0 U1546 ( .I0(n1576), .I1(rw_C1_M[1]), .S(n1575), .ZN(n1577) );
  HVT_OA21HSV2 U1549 ( .A1(n1669), .A2(n1676), .B(1'b0), .Z(n1073) );
  LVT_NAND3HSV2 U1556 ( .A1(n148), .A2(n3039), .A3(n449), .ZN(n447) );
  LVT_INOR2HSV1 U1559 ( .A1(n801), .B1(n3047), .ZN(n697) );
  LVT_OAI211HSV1 U1560 ( .A1(n656), .A2(n657), .B(n664), .C(n1865), .ZN(n659)
         );
  HVT_OAI22HSV0 U1561 ( .A1(n438), .A2(n2560), .B1(n439), .B2(n3091), .ZN(
        n1040) );
  HVT_AOI211HSV0 U1563 ( .A1(n3099), .A2(n3074), .B(n456), .C(n691), .ZN(n689)
         );
  HVT_AOI211HSV0 U1564 ( .A1(n3058), .A2(n1804), .B(n3044), .C(n1802), .ZN(
        n587) );
  LVT_INOR2HSV1 U1565 ( .A1(n552), .B1(n550), .ZN(n551) );
  LVT_INOR2HSV1 U1566 ( .A1(n654), .B1(n652), .ZN(n653) );
  LVT_NOR2HSV2 U1567 ( .A1(n701), .A2(n713), .ZN(n700) );
  LVT_MUX2NHSV1 U1585 ( .I0(n1466), .I1(n3098), .S(n155), .ZN(n1173) );
  LVT_MUX2NHSV1 U1587 ( .I0(n3067), .I1(n1484), .S(n659), .ZN(n1152) );
  LVT_AND3HSV2 U1588 ( .A1(n655), .A2(n1865), .A3(n657), .Z(n1484) );
  LVT_NAND2HSV2 U1589 ( .A1(n1812), .A2(n1811), .ZN(n575) );
  LVT_INOR2HSV1 U1590 ( .A1(n513), .B1(n577), .ZN(n1812) );
  LVT_MUX2NHSV1 U1591 ( .I0(n1580), .I1(n2452), .S(n1579), .ZN(n1175) );
  LVT_NAND2HSV2 U1614 ( .A1(n528), .A2(n529), .ZN(n1076) );
  HVT_AOI211HSV0 U1615 ( .A1(n3069), .A2(n3075), .B(n527), .C(n536), .ZN(n528)
         );
  LVT_NAND2HSV2 U1618 ( .A1(n736), .A2(n737), .ZN(n1190) );
  HVT_AOI211HSV0 U1619 ( .A1(n522), .A2(n500), .B(n501), .C(n424), .ZN(n736)
         );
  HVT_OAI211HSV0 U1621 ( .A1(n1674), .A2(n3063), .B(n1672), .C(n1671), .ZN(
        n1675) );
  LVT_NAND2HSV2 U1622 ( .A1(n630), .A2(n631), .ZN(n1126) );
  LVT_INOR2HSV1 U1623 ( .A1(n650), .B1(n160), .ZN(n649) );
  HVT_OAI22HSV0 U1625 ( .A1(n438), .A2(n2466), .B1(n439), .B2(n3087), .ZN(
        n1047) );
  HVT_OAI22HSV0 U1626 ( .A1(n438), .A2(n2467), .B1(n439), .B2(n3094), .ZN(
        n1043) );
  HVT_OAI22HSV0 U1627 ( .A1(n438), .A2(n2556), .B1(n439), .B2(n3086), .ZN(
        n1041) );
  LVT_AND3HSV2 U1630 ( .A1(n1849), .A2(n1818), .A3(n1817), .Z(n539) );
  HVT_OAI22HSV0 U1632 ( .A1(n438), .A2(n2438), .B1(n3092), .B2(n439), .ZN(
        n1052) );
  HVT_OAI22HSV0 U1633 ( .A1(n438), .A2(n2462), .B1(n3089), .B2(n439), .ZN(
        n1051) );
  HVT_OAI22HSV0 U1634 ( .A1(n438), .A2(n2461), .B1(n3095), .B2(n439), .ZN(
        n1050) );
  HVT_OAI22HSV0 U1635 ( .A1(n438), .A2(n1294), .B1(n3093), .B2(n439), .ZN(
        n1042) );
  HVT_OAI22HSV0 U1636 ( .A1(n438), .A2(n2459), .B1(n3085), .B2(n439), .ZN(
        n1037) );
  LVT_OAI211HSV1 U1640 ( .A1(n592), .A2(n591), .B(n1664), .C(n1663), .ZN(n1802) );
  LVT_OAI221HSV1 U1643 ( .A1(en_C2_P2), .A2(n555), .B1(n570), .B2(n561), .C(
        n1855), .ZN(n1105) );
  LVT_OAI221HSV1 U1645 ( .A1(en_C1_P1), .A2(n657), .B1(n672), .B2(n663), .C(
        n1866), .ZN(n1155) );
  LVT_INOR3HSV2 U1647 ( .A1(debugRwToMem[1]), .B1(debugRwToMem[0]), .B2(reset), 
        .ZN(n713) );
  LVT_AO32HSV1 U1648 ( .A1(n157), .A2(n712), .A3(n707), .B1(n1018), .B2(
        mb_chipSelect), .Z(n1211) );
  LVT_OA221HSV2 U1652 ( .A1(n553), .A2(n161), .B1(n554), .B2(n555), .C(C1_N80), 
        .Z(n550) );
  LVT_OA221HSV2 U1653 ( .A1(n655), .A2(n160), .B1(n656), .B2(n657), .C(C1_N80), 
        .Z(n652) );
  LVT_NAND2HSV2 U1655 ( .A1(n569), .A2(stateP2[0]), .ZN(n561) );
  HVT_MOAI22HSV0 U1656 ( .A1(n547), .A2(n3092), .B1(ins_code2_proc2[0]), .B2(
        n547), .ZN(n1093) );
  LVT_NAND2HSV2 U1658 ( .A1(n671), .A2(stateP1[0]), .ZN(n663) );
  LVT_OAI211HSV1 U1659 ( .A1(n554), .A2(n555), .B(n1693), .C(n1692), .ZN(n1694) );
  LVT_INOR2HSV1 U1660 ( .A1(n548), .B1(n161), .ZN(n547) );
  LVT_AOI211HSV1 U1661 ( .A1(n641), .A2(n3055), .B(reset), .C(n2570), .ZN(n640) );
  LVT_NOR2HSV2 U1662 ( .A1(debugRwToMem[1]), .A2(reset), .ZN(n699) );
  LVT_MUX2NHSV1 U1663 ( .I0(n3066), .I1(n1486), .S(n659), .ZN(n1153) );
  LVT_AND4HSV2 U1664 ( .A1(n553), .A2(C1_N80), .A3(n1696), .A4(n555), .Z(n1698) );
  LVT_MUX2NHSV1 U1665 ( .I0(n1455), .I1(n1457), .S(debugDelay[5]), .ZN(n1178)
         );
  LVT_MUX2NHSV1 U1666 ( .I0(n1460), .I1(n1461), .S(debugDelay[6]), .ZN(n1177)
         );
  LVT_MUX2NHSV1 U1667 ( .I0(n159), .I1(n2474), .S(n700), .ZN(n1174) );
  LVT_MUX2NHSV1 U1668 ( .I0(n1445), .I1(n1444), .S(debugDelay[3]), .ZN(n1180)
         );
  LVT_AOI211HSV1 U1674 ( .A1(n2411), .A2(n3068), .B(n729), .C(n2512), .ZN(
        n1714) );
  HVT_NAND2HSV0 U1675 ( .A1(n639), .A2(C1_N80), .ZN(n729) );
  HVT_OAI211HSV0 U1677 ( .A1(n1674), .A2(n3061), .B(n1655), .C(n1654), .ZN(
        n1656) );
  LVT_IOA21HSV2 U1680 ( .A1(n1359), .A2(en_C1_P1), .B(n1790), .ZN(n1156) );
  LVT_INOR2HSV1 U1684 ( .A1(n673), .B1(reset), .ZN(n671) );
  LVT_NOR2HSV2 U1686 ( .A1(n561), .A2(ins_code2_proc2[23]), .ZN(n556) );
  LVT_INOR2HSV1 U1687 ( .A1(n571), .B1(reset), .ZN(n569) );
  LVT_NOR2HSV2 U1688 ( .A1(n663), .A2(ins_code1_proc1[23]), .ZN(n658) );
  LVT_IOA22HSV1 U1692 ( .B1(n700), .B2(n708), .A1(debugRwToMem[1]), .A2(n700), 
        .ZN(n1185) );
  LVT_INOR4HSV2 U1693 ( .A1(n1871), .B1(mb_stall), .B2(n709), .B3(n710), .ZN(
        n708) );
  LVT_INOR4HSV2 U1697 ( .A1(n417), .B1(n418), .B2(n3046), .B3(reset), .ZN(n416) );
  LVT_OAI221HSV1 U1698 ( .A1(n571), .A2(reset), .B1(n565), .B2(n555), .C(n1685), .ZN(n1686) );
  LVT_OAI221HSV1 U1699 ( .A1(n673), .A2(reset), .B1(n667), .B2(n657), .C(n1475), .ZN(n1476) );
  LVT_AOI21HSV2 U1713 ( .A1(n542), .A2(n543), .B(reset), .ZN(n1077) );
  HVT_MUX2NHSV0 U1716 ( .I0(addr_P1_C1[0]), .I1(ins_code1_proc1[0]), .S(n649), 
        .ZN(n1485) );
  HVT_MUX2NHSV0 U1717 ( .I0(addr_P1_C1[1]), .I1(ins_code1_proc1[1]), .S(n649), 
        .ZN(n1524) );
  HVT_MUX2NHSV0 U1718 ( .I0(addr_P1_C1[2]), .I1(ins_code1_proc1[2]), .S(n649), 
        .ZN(n1523) );
  HVT_MUX2NHSV0 U1719 ( .I0(addr_P1_C1[3]), .I1(ins_code1_proc1[3]), .S(n649), 
        .ZN(n1488) );
  HVT_MUX2NHSV0 U1720 ( .I0(addr_P1_C1[4]), .I1(ins_code1_proc1[4]), .S(n649), 
        .ZN(n1528) );
  HVT_MUX2NHSV0 U1721 ( .I0(addr_P1_C1[5]), .I1(ins_code1_proc1[5]), .S(n649), 
        .ZN(n1527) );
  HVT_MUX2NHSV0 U1722 ( .I0(addr_P1_C1[6]), .I1(ins_code1_proc1[6]), .S(n649), 
        .ZN(n1526) );
  HVT_MUX2NHSV0 U1723 ( .I0(addr_P1_C1[9]), .I1(ins_code1_proc1[9]), .S(n649), 
        .ZN(n1530) );
  HVT_MUX2NHSV0 U1724 ( .I0(addr_P1_C1[10]), .I1(ins_code1_proc1[10]), .S(n649), .ZN(n1529) );
  HVT_MUX2NHSV0 U1725 ( .I0(addr_P1_C1[12]), .I1(ins_code1_proc1[12]), .S(n649), .ZN(n1535) );
  HVT_MUX2NHSV0 U1726 ( .I0(addr_P1_C1[13]), .I1(ins_code1_proc1[13]), .S(n649), .ZN(n1534) );
  HVT_MUX2NHSV0 U1727 ( .I0(addr_P1_C1[14]), .I1(ins_code1_proc1[14]), .S(n649), .ZN(n1533) );
  HVT_MUX2NHSV0 U1728 ( .I0(addr_P1_C1[15]), .I1(ins_code1_proc1[15]), .S(n649), .ZN(n1525) );
  HVT_MUX2NHSV0 U1729 ( .I0(addr_P2_C2[1]), .I1(ins_code2_proc2[1]), .S(n547), 
        .ZN(n1405) );
  HVT_MUX2NHSV0 U1730 ( .I0(addr_P2_C2[2]), .I1(ins_code2_proc2[2]), .S(n547), 
        .ZN(n1407) );
  HVT_MUX2NHSV0 U1731 ( .I0(n1290), .I1(ins_code2_proc2[3]), .S(n547), .ZN(
        n1427) );
  HVT_MUX2NHSV0 U1732 ( .I0(addr_P2_C2[5]), .I1(ins_code2_proc2[5]), .S(n547), 
        .ZN(n1425) );
  HVT_MUX2NHSV0 U1733 ( .I0(addr_P2_C2[6]), .I1(ins_code2_proc2[6]), .S(n547), 
        .ZN(n1424) );
  HVT_MUX2NHSV0 U1734 ( .I0(addr_P2_C2[7]), .I1(ins_code2_proc2[7]), .S(n547), 
        .ZN(n1419) );
  HVT_MUX2NHSV0 U1735 ( .I0(addr_P2_C2[8]), .I1(ins_code2_proc2[8]), .S(n547), 
        .ZN(n1418) );
  HVT_MUX2NHSV0 U1736 ( .I0(addr_P2_C2[9]), .I1(ins_code2_proc2[9]), .S(n547), 
        .ZN(n1417) );
  HVT_MUX2NHSV0 U1737 ( .I0(addr_P2_C2[11]), .I1(ins_code2_proc2[11]), .S(n547), .ZN(n1411) );
  HVT_MUX2NHSV0 U1738 ( .I0(addr_P2_C2[13]), .I1(ins_code2_proc2[13]), .S(n547), .ZN(n1409) );
  HVT_MUX2NHSV0 U1739 ( .I0(addr_P2_C2[14]), .I1(ins_code2_proc2[14]), .S(n547), .ZN(n1408) );
  HVT_MUX2NHSV0 U1740 ( .I0(addr_P2_C2[15]), .I1(ins_code2_proc2[15]), .S(n547), .ZN(n1404) );
  HVT_MUX2NHSV0 U1741 ( .I0(addr_P1_C1[7]), .I1(ins_code1_proc1[7]), .S(n649), 
        .ZN(n1532) );
  LVT_MUX2NHSV1 U1742 ( .I0(n1432), .I1(n1452), .S(debugDelay[0]), .ZN(n1433)
         );
  LVT_AOI21HSV2 U1743 ( .A1(en_M_C1), .A2(n3045), .B(n604), .ZN(n719) );
  LVT_OA21HSV2 U1763 ( .A1(n148), .A2(n414), .B(1'b0), .Z(n1054) );
  LVT_INAND2HSV2 U1766 ( .A1(reset), .B1(n1569), .ZN(n1517) );
  HVT_MUX2NHSV0 U1769 ( .I0(addr_P2_C2[4]), .I1(ins_code2_proc2[4]), .S(n547), 
        .ZN(n1426) );
  HVT_AOI31HSV0 U1773 ( .A1(n3078), .A2(n3077), .A3(n3070), .B(n527), .ZN(n510) );
  HVT_AND4HSV1 U1779 ( .A1(n463), .A2(msg_C1_C2), .A3(C1_N80), .A4(n3050), .Z(
        n1654) );
  HVT_OAI211HSV0 U1780 ( .A1(n1543), .A2(n1553), .B(n3050), .C(n1542), .ZN(
        n1544) );
  HVT_MUX2NHSV0 U1787 ( .I0(addr_P1_C1[8]), .I1(ins_code1_proc1[8]), .S(n649), 
        .ZN(n1531) );
  LVT_AO22HSV1 U1788 ( .A1(n1659), .A2(addr_P1_C1[8]), .B1(addr_C1_C2[8]), 
        .B2(n1658), .Z(n1063) );
  HVT_MUX2NHSV0 U1791 ( .I0(addr_P1_C1[11]), .I1(ins_code1_proc1[11]), .S(n649), .ZN(n1536) );
  HVT_OAI21HSV0 U1796 ( .A1(n1662), .A2(n1635), .B(n1634), .ZN(n1636) );
  LVT_OAI222HSV0 U1816 ( .A1(n1916), .A2(n435), .B1(n1277), .B2(n436), .C1(
        n437), .C2(n2477), .ZN(n1033) );
  LVT_OAI222HSV0 U1817 ( .A1(n1916), .A2(n695), .B1(n1277), .B2(n696), .C1(
        n697), .C2(n2426), .ZN(n1169) );
  LVT_OAI222HSV0 U1818 ( .A1(n3086), .A2(n695), .B1(n2563), .B2(n696), .C1(
        n697), .C2(n2446), .ZN(n1161) );
  HVT_OAI222HSV0 U1819 ( .A1(n3086), .A2(n435), .B1(n2563), .B2(n436), .C1(
        n437), .C2(n2472), .ZN(n1025) );
  LVT_OAI222HSV0 U1822 ( .A1(n2562), .A2(n695), .B1(n2533), .B2(n696), .C1(
        n697), .C2(n2445), .ZN(n1159) );
  LVT_OAI22HSV0 U1823 ( .A1(n438), .A2(n2412), .B1(n2562), .B2(n439), .ZN(
        n1039) );
  HVT_OAI222HSV0 U1824 ( .A1(n2562), .A2(n435), .B1(n2533), .B2(n436), .C1(
        n437), .C2(n2505), .ZN(n1023) );
  LVT_OAI21HSV4 U1826 ( .A1(n1250), .A2(n2011), .B(n1818), .ZN(n1658) );
  LVT_OR4HSV2 U1828 ( .A1(n1228), .A2(n2011), .A3(n3045), .A4(n1785), .Z(n1788) );
  HVT_OAI222HSV0 U1832 ( .A1(n3090), .A2(n435), .B1(n3079), .B2(n436), .C1(
        n437), .C2(n2469), .ZN(n1029) );
  LVT_OAI222HSV0 U1833 ( .A1(n3090), .A2(n695), .B1(n3079), .B2(n696), .C1(
        n697), .C2(n2442), .ZN(n1165) );
  HVT_OAI222HSV0 U1837 ( .A1(n3096), .A2(n435), .B1(n3081), .B2(n436), .C1(
        n437), .C2(n2479), .ZN(n1030) );
  LVT_OAI222HSV0 U1838 ( .A1(n3096), .A2(n695), .B1(n3081), .B2(n696), .C1(
        n697), .C2(n2443), .ZN(n1166) );
  LVT_OAI222HSV0 U1839 ( .A1(n2395), .A2(n695), .B1(n2535), .B2(n696), .C1(
        n697), .C2(n2449), .ZN(n1158) );
  LVT_OAI22HSV0 U1840 ( .A1(n438), .A2(n2403), .B1(n2395), .B2(n439), .ZN(
        n1038) );
  HVT_OAI222HSV0 U1841 ( .A1(n2395), .A2(n435), .B1(n2535), .B2(n436), .C1(
        n437), .C2(n2504), .ZN(n1022) );
  LVT_OAI222HSV0 U1845 ( .A1(n3088), .A2(n695), .B1(n3080), .B2(n696), .C1(
        n697), .C2(n2440), .ZN(n1164) );
  HVT_OAI222HSV0 U1848 ( .A1(n3097), .A2(n435), .B1(n2546), .B2(n436), .C1(
        n437), .C2(n2478), .ZN(n1032) );
  LVT_OAI222HSV0 U1849 ( .A1(n3097), .A2(n695), .B1(n2546), .B2(n696), .C1(
        n697), .C2(n2444), .ZN(n1168) );
  HVT_MUX2NHSV0 U1850 ( .I0(addr_P2_C2[12]), .I1(ins_code2_proc2[12]), .S(n547), .ZN(n1410) );
  HVT_MUX2NHSV0 U1855 ( .I0(addr_P2_C2[10]), .I1(ins_code2_proc2[10]), .S(n547), .ZN(n1416) );
  LVT_OAI22HSV2 U1856 ( .A1(n438), .A2(n2460), .B1(n1916), .B2(n439), .ZN(
        n1049) );
  HVT_AND2HSV2 U1857 ( .A1(n431), .A2(n1737), .Z(n1738) );
  LVT_OAI22HSV2 U1861 ( .A1(n438), .A2(n2558), .B1(n3090), .B2(n439), .ZN(
        n1045) );
  LVT_OAI22HSV2 U1862 ( .A1(n438), .A2(n2559), .B1(n3096), .B2(n439), .ZN(
        n1046) );
  LVT_OAI22HSV2 U1863 ( .A1(n438), .A2(n2458), .B1(n3088), .B2(n439), .ZN(
        n1044) );
  LVT_OAI22HSV2 U1865 ( .A1(n438), .A2(n2457), .B1(n3097), .B2(n439), .ZN(
        n1048) );
  LVT_CLKNHSV2 U1868 ( .I(n1404), .ZN(n1078) );
  LVT_CLKNHSV2 U1869 ( .I(n1405), .ZN(n1092) );
  LVT_CLKNHSV2 U1870 ( .I(n1407), .ZN(n1091) );
  LVT_CLKNHSV2 U1871 ( .I(n1408), .ZN(n1079) );
  LVT_CLKNHSV2 U1872 ( .I(n1409), .ZN(n1080) );
  LVT_CLKNHSV2 U1873 ( .I(n1410), .ZN(n1081) );
  LVT_CLKNHSV2 U1874 ( .I(n1411), .ZN(n1082) );
  LVT_CLKNHSV2 U1876 ( .I(n1416), .ZN(n1083) );
  LVT_CLKNHSV2 U1877 ( .I(n1417), .ZN(n1084) );
  LVT_CLKNHSV2 U1878 ( .I(n1418), .ZN(n1085) );
  LVT_CLKNHSV2 U1879 ( .I(n1419), .ZN(n1086) );
  LVT_CLKNHSV2 U1881 ( .I(n1424), .ZN(n1087) );
  LVT_CLKNHSV2 U1882 ( .I(n1425), .ZN(n1088) );
  LVT_CLKNHSV2 U1883 ( .I(n1426), .ZN(n1089) );
  LVT_CLKNHSV2 U1884 ( .I(n1427), .ZN(n1090) );
  LVT_OAI21HSV2 U1892 ( .A1(n159), .A2(n1434), .B(C1_N80), .ZN(n701) );
  LVT_CLKNHSV2 U1893 ( .I(n699), .ZN(n1432) );
  LVT_INAND2HSV2 U1894 ( .A1(reset), .B1(n1432), .ZN(n1452) );
  LVT_CLKNHSV2 U1895 ( .I(n701), .ZN(n1579) );
  LVT_INAND2HSV2 U1896 ( .A1(n1433), .B1(n1579), .ZN(n1183) );
  LVT_INAND2HSV2 U1897 ( .A1(n159), .B1(n1434), .ZN(n1464) );
  LVT_CLKNHSV2 U1898 ( .I(n1464), .ZN(n1448) );
  LVT_CLKNHSV2 U1901 ( .I(n1452), .ZN(n1871) );
  LVT_AO22HSV0 U1902 ( .A1(n1448), .A2(n1438), .B1(debugDelay[1]), .B2(n1871), 
        .Z(n1182) );
  LVT_AO221HSV0 U1905 ( .A1(n699), .A2(n1441), .B1(n1871), .B2(debugDelay[2]), 
        .C(n701), .Z(n1181) );
  LVT_INAND2HSV2 U1906 ( .A1(n1442), .B1(n1448), .ZN(n1445) );
  LVT_OAI21HSV2 U1908 ( .A1(n2451), .A2(n1464), .B(n1452), .ZN(n1446) );
  LVT_CLKNHSV2 U1909 ( .I(n1446), .ZN(n1444) );
  LVT_IAO21HSV0 U1911 ( .A1(n1464), .A2(n2485), .B(n1446), .ZN(n1450) );
  LVT_INAND2HSV2 U1913 ( .A1(n1451), .B1(n1448), .ZN(n1455) );
  LVT_OAI21HSV2 U1914 ( .A1(n1450), .A2(n2434), .B(n1455), .ZN(n1179) );
  LVT_OAI21HSV2 U1916 ( .A1(n2435), .A2(n1464), .B(n1452), .ZN(n1454) );
  LVT_CLKNHSV2 U1917 ( .I(n1454), .ZN(n1457) );
  LVT_CLKNHSV2 U1918 ( .I(n1455), .ZN(n1456) );
  LVT_INAND2HSV2 U1919 ( .A1(debugDelay[5]), .B1(n1456), .ZN(n1460) );
  LVT_OAI21HSV2 U1921 ( .A1(n1464), .A2(n2501), .B(n1457), .ZN(n1459) );
  LVT_CLKNHSV2 U1922 ( .I(n1459), .ZN(n1461) );
  LVT_OAI32HSV2 U1925 ( .A1(n1464), .A2(n2484), .A3(1'b1), .B1(n1461), .B2(
        1'b1), .ZN(n1176) );
  LVT_INAND2HSV2 U1927 ( .A1(mb_stall), .B1(n713), .ZN(n1588) );
  LVT_INAND2HSV2 U1928 ( .A1(n701), .B1(n1588), .ZN(n698) );
  LVT_INAND2HSV2 U1930 ( .A1(n2463), .B1(n699), .ZN(n1466) );
  LVT_CLKNHSV2 U1932 ( .I(n698), .ZN(n155) );
  LVT_OAI222HSV2 U1944 ( .A1(n695), .A2(n3092), .B1(n696), .B2(n3082), .C1(
        n697), .C2(n2437), .ZN(n1172) );
  LVT_INAND2HSV2 U1945 ( .A1(stateP1[0]), .B1(n671), .ZN(n1478) );
  LVT_INAND2HSV2 U1946 ( .A1(n1478), .B1(stateP1[1]), .ZN(n657) );
  LVT_CLKNHSV2 U1947 ( .I(n657), .ZN(n1471) );
  LVT_INAND2HSV2 U1948 ( .A1(n1471), .B1(n663), .ZN(n654) );
  LVT_OAI21HSV2 U1950 ( .A1(n2591), .A2(n663), .B(n657), .ZN(n1474) );
  LVT_CLKNHSV2 U1951 ( .I(n654), .ZN(n1473) );
  LVT_IAO22HSV1 U1953 ( .B1(ins_code1_proc1[22]), .B2(n1474), .A1(n1473), .A2(
        n2588), .ZN(n1475) );
  LVT_CLKNHSV2 U1954 ( .I(n1476), .ZN(n1866) );
  LVT_OAI31HSV2 U1955 ( .A1(n2590), .A2(n663), .A3(n2592), .B(n1866), .ZN(
        n1480) );
  LVT_CLKNHSV2 U1956 ( .I(n1478), .ZN(n1479) );
  LVT_INAND2HSV2 U1957 ( .A1(stateP1[1]), .B1(n1479), .ZN(n1481) );
  LVT_INAND2HSV2 U1958 ( .A1(n1480), .B1(n1481), .ZN(n1154) );
  LVT_CLKNHSV2 U1960 ( .I(n1481), .ZN(n1482) );
  LVT_INAND2HSV2 U1961 ( .A1(n1482), .B1(C1_N80), .ZN(n1483) );
  LVT_CLKNHSV2 U1962 ( .I(n1483), .ZN(n1865) );
  LVT_CLKNHSV2 U1963 ( .I(n1485), .ZN(n1143) );
  LVT_INAND2HSV2 U1965 ( .A1(n663), .B1(n666), .ZN(n1486) );
  LVT_CLKNHSV2 U1966 ( .I(n1488), .ZN(n1140) );
  LVT_CLKNHSV2 U1985 ( .I(n1517), .ZN(n1521) );
  LVT_INAND2HSV2 U1986 ( .A1(n1624), .B1(n1521), .ZN(n1539) );
  LVT_INAND2HSV2 U1988 ( .A1(n3056), .B1(n1521), .ZN(n1518) );
  LVT_CLKNHSV2 U1989 ( .I(n1518), .ZN(n1538) );
  LVT_OAI31HSV2 U1995 ( .A1(n3049), .A2(n3041), .A3(n1635), .B(n1521), .ZN(
        n1537) );
  LVT_OAI222HSV2 U1996 ( .A1(n2540), .A2(n1539), .B1(n1538), .B2(n2422), .C1(
        n2581), .C2(n1537), .ZN(n1119) );
  LVT_CLKNHSV2 U1998 ( .I(n1523), .ZN(n1141) );
  LVT_OAI222HSV2 U2001 ( .A1(n2539), .A2(n1539), .B1(n1538), .B2(n2423), .C1(
        n2549), .C2(n1537), .ZN(n1120) );
  LVT_CLKNHSV2 U2002 ( .I(n1524), .ZN(n1142) );
  LVT_OAI222HSV2 U2006 ( .A1(n2555), .A2(n1539), .B1(n1538), .B2(n2424), .C1(
        n2551), .C2(n1537), .ZN(n1121) );
  LVT_OAI32HSV2 U2007 ( .A1(n3032), .A2(n147), .A3(reset), .B1(n447), .B2(
        n2483), .ZN(n1053) );
  LVT_OAI222HSV2 U2011 ( .A1(n3057), .A2(n1539), .B1(n1538), .B2(n2415), .C1(
        n3059), .C2(n1537), .ZN(n1122) );
  LVT_CLKNHSV2 U2012 ( .I(n1525), .ZN(n1128) );
  LVT_OAI222HSV2 U2015 ( .A1(n2580), .A2(n1539), .B1(n1538), .B2(n2425), .C1(
        n2577), .C2(n1537), .ZN(n1207) );
  LVT_CLKNHSV2 U2016 ( .I(n1526), .ZN(n1137) );
  LVT_OAI222HSV2 U2018 ( .A1(n2538), .A2(n1539), .B1(n1538), .B2(n2432), .C1(
        n2557), .C2(n1537), .ZN(n1116) );
  LVT_CLKNHSV2 U2019 ( .I(n1527), .ZN(n1138) );
  LVT_OAI222HSV2 U2021 ( .A1(n2542), .A2(n1539), .B1(n1538), .B2(n2433), .C1(
        n2550), .C2(n1537), .ZN(n1117) );
  LVT_CLKNHSV2 U2022 ( .I(n1528), .ZN(n1139) );
  LVT_OAI222HSV2 U2025 ( .A1(n2579), .A2(n1539), .B1(n1538), .B2(n2421), .C1(
        n2578), .C2(n1537), .ZN(n1118) );
  LVT_CLKNHSV2 U2026 ( .I(n1529), .ZN(n1133) );
  LVT_OAI222HSV2 U2029 ( .A1(n2524), .A2(n1539), .B1(n1538), .B2(n2429), .C1(
        n2529), .C2(n1537), .ZN(n1112) );
  LVT_CLKNHSV2 U2030 ( .I(n1530), .ZN(n1134) );
  LVT_OAI222HSV2 U2033 ( .A1(n2521), .A2(n1539), .B1(n1538), .B2(n2430), .C1(
        n2531), .C2(n1537), .ZN(n1113) );
  LVT_CLKNHSV2 U2034 ( .I(n1531), .ZN(n1135) );
  LVT_OAI222HSV2 U2037 ( .A1(n2541), .A2(n1539), .B1(n1538), .B2(n2420), .C1(
        n2530), .C2(n1537), .ZN(n1114) );
  LVT_CLKNHSV2 U2038 ( .I(n1532), .ZN(n1136) );
  LVT_OAI222HSV2 U2041 ( .A1(n2522), .A2(n1539), .B1(n1538), .B2(n2431), .C1(
        n2514), .C2(n1537), .ZN(n1115) );
  LVT_CLKNHSV2 U2042 ( .I(n1533), .ZN(n1129) );
  LVT_OAI222HSV2 U2045 ( .A1(n2545), .A2(n1539), .B1(n1538), .B2(n2417), .C1(
        n2509), .C2(n1537), .ZN(n1108) );
  LVT_CLKNHSV2 U2046 ( .I(n1534), .ZN(n1130) );
  LVT_OAI222HSV2 U2049 ( .A1(n1281), .A2(n1539), .B1(n1538), .B2(n2418), .C1(
        n2575), .C2(n1537), .ZN(n1109) );
  LVT_CLKNHSV2 U2050 ( .I(n1535), .ZN(n1131) );
  LVT_OAI222HSV2 U2053 ( .A1(n1297), .A2(n1539), .B1(n1538), .B2(n2419), .C1(
        n2574), .C2(n1537), .ZN(n1110) );
  LVT_CLKNHSV2 U2054 ( .I(n1536), .ZN(n1132) );
  LVT_OAI222HSV2 U2056 ( .A1(n1279), .A2(n1539), .B1(n1538), .B2(n2428), .C1(
        n2576), .C2(n1537), .ZN(n1111) );
  LVT_CLKNHSV2 U2060 ( .I(n604), .ZN(n1542) );
  LVT_INAND2HSV2 U2061 ( .A1(n3065), .B1(n1544), .ZN(n1547) );
  LVT_CLKNHSV2 U2062 ( .I(C1_N80), .ZN(n1840) );
  LVT_INAND2HSV2 U2063 ( .A1(reset), .B1(n3056), .ZN(n1787) );
  LVT_CLKNHSV2 U2064 ( .I(n1787), .ZN(n1676) );
  LVT_CLKNHSV2 U2065 ( .I(n1544), .ZN(n1545) );
  LVT_OAI21HSV2 U2066 ( .A1(n1676), .A2(n1545), .B(C1_stall), .ZN(n1546) );
  LVT_OAI31HSV2 U2067 ( .A1(n1547), .A2(n600), .A3(n1840), .B(n1546), .ZN(
        n1124) );
  LVT_AO221HSV0 U2073 ( .A1(n3054), .A2(n3065), .B1(n3064), .B2(n3062), .C(
        n1556), .Z(n1792) );
  LVT_OR3HSV0 U2075 ( .A1(n3041), .A2(n1792), .A3(n3040), .Z(n1561) );
  LVT_INAND2HSV2 U2076 ( .A1(n1564), .B1(n1563), .ZN(n1125) );
  LVT_CLKNHSV2 U2079 ( .I(reset), .ZN(n1818) );
  LVT_CLKAND2HSV2 U2080 ( .A1(n1568), .A2(n1818), .Z(n1127) );
  LVT_CLKNHSV2 U2081 ( .I(n719), .ZN(n151) );
  LVT_CLKNHSV2 U2082 ( .I(n1570), .ZN(n1575) );
  LVT_OAI21HSV2 U2083 ( .A1(n1676), .A2(n1575), .B(rw_C1_M[0]), .ZN(n1571) );
  LVT_OAI21HSV2 U2084 ( .A1(n1840), .A2(n1624), .B(n1571), .ZN(n1123) );
  LVT_OR4HSV0 U2086 ( .A1(reset), .A2(n3051), .A3(n716), .A4(n3045), .Z(n1576)
         );
  LVT_CLKNHSV2 U2087 ( .I(n1577), .ZN(n1186) );
  LVT_INAND2HSV2 U2089 ( .A1(n159), .B1(n2463), .ZN(n1580) );
  LVT_OAI21HSV2 U2094 ( .A1(n3098), .A2(n1849), .B(C1_N80), .ZN(n577) );
  LVT_INAND2HSV2 U2098 ( .A1(n577), .B1(n1780), .ZN(n424) );
  LVT_CLKNHSV2 U2099 ( .I(n1585), .ZN(n1857) );
  LVT_INAND2HSV2 U2100 ( .A1(n420), .B1(n1818), .ZN(n1586) );
  LVT_CLKNHSV2 U2101 ( .I(n1586), .ZN(n414) );
  LVT_OAI21HSV2 U2102 ( .A1(n1857), .A2(n414), .B(rw_C2_M[0]), .ZN(n1587) );
  LVT_CLKNHSV2 U2104 ( .I(n1588), .ZN(n1870) );
  LVT_AO22HSV0 U2109 ( .A1(n1870), .A2(n1592), .B1(debugRwToMem[0]), .B2(n700), 
        .Z(n1184) );
  LVT_INAND2HSV2 U2115 ( .A1(reset), .B1(n2407), .ZN(n873) );
  LVT_OR3HSV0 U2116 ( .A1(reset), .A2(n3056), .A3(n3048), .Z(n1627) );
  LVT_CLKNHSV2 U2117 ( .I(n1627), .ZN(n874) );
  LVT_OAI222HSV2 U2119 ( .A1(n873), .A2(n3057), .B1(n872), .B2(n3059), .C1(
        n874), .C2(n2500), .ZN(n1206) );
  LVT_CLKNHSV2 U2136 ( .I(n1658), .ZN(n1634) );
  LVT_CLKNHSV2 U2137 ( .I(n1636), .ZN(n1659) );
  LVT_AO22HSV0 U2138 ( .A1(n1659), .A2(addr_P1_C1[7]), .B1(addr_C1_C2[7]), 
        .B2(n1658), .Z(n1064) );
  LVT_AO22HSV0 U2139 ( .A1(n1659), .A2(addr_P1_C1[10]), .B1(addr_C1_C2[10]), 
        .B2(n1658), .Z(n1061) );
  LVT_OAI21HSV2 U2142 ( .A1(reset), .A2(n1657), .B(n1656), .ZN(n1055) );
  LVT_AO22HSV0 U2143 ( .A1(n1659), .A2(addr_P1_C1[14]), .B1(addr_C1_C2[14]), 
        .B2(n1658), .Z(n1057) );
  LVT_CLKAND2HSV2 U2144 ( .A1(C1_N80), .A2(n683), .Z(n1663) );
  LVT_CLKNHSV2 U2145 ( .I(n1802), .ZN(n1669) );
  LVT_CLKAND2HSV2 U2147 ( .A1(n3052), .A2(n1669), .Z(n1671) );
  LVT_CLKNHSV2 U2148 ( .I(n1675), .ZN(n1678) );
  LVT_OAI21HSV2 U2149 ( .A1(n1676), .A2(n1678), .B(wm_C1_C2), .ZN(n1677) );
  LVT_OAI31HSV2 U2150 ( .A1(n1679), .A2(reset), .A3(n1678), .B(n1677), .ZN(
        n1072) );
  LVT_CLKNHSV2 U2152 ( .I(n569), .ZN(n1687) );
  LVT_OR3HSV0 U2153 ( .A1(n2465), .A2(n1687), .A3(stateP2[0]), .Z(n555) );
  LVT_CLKNHSV2 U2154 ( .I(n555), .ZN(n1681) );
  LVT_INAND2HSV2 U2155 ( .A1(n1681), .B1(n561), .ZN(n552) );
  LVT_OAI21HSV2 U2157 ( .A1(n2586), .A2(n561), .B(n555), .ZN(n1684) );
  LVT_CLKNHSV2 U2158 ( .I(n552), .ZN(n1683) );
  LVT_IAO22HSV1 U2160 ( .B1(ins_code2_proc2[22]), .B2(n1684), .A1(n1683), .A2(
        n2582), .ZN(n1685) );
  LVT_CLKNHSV2 U2161 ( .I(n1686), .ZN(n1855) );
  LVT_OR3HSV0 U2162 ( .A1(stateP2[0]), .A2(n1687), .A3(stateP2[1]), .Z(n1696)
         );
  LVT_CLKAND2HSV2 U2163 ( .A1(n1855), .A2(n1696), .Z(n1688) );
  LVT_OAI31HSV2 U2164 ( .A1(n2584), .A2(n561), .A3(n2587), .B(n1688), .ZN(
        n1104) );
  LVT_CLKNHSV2 U2168 ( .I(n561), .ZN(n1691) );
  LVT_INAND2HSV2 U2169 ( .A1(n2585), .B1(n1691), .ZN(n1695) );
  LVT_OAI31HSV2 U2171 ( .A1(n2583), .A2(n564), .A3(n560), .B(n556), .ZN(n1693)
         );
  LVT_CLKAND2HSV2 U2172 ( .A1(C1_N80), .A2(n1696), .Z(n1692) );
  LVT_CLKNHSV2 U2173 ( .I(n1694), .ZN(n1697) );
  LVT_CLKNHSV2 U2174 ( .I(n1708), .ZN(n1715) );
  LVT_OAI21HSV2 U2176 ( .A1(n3056), .A2(n1715), .B(allowRead_C1_C2), .ZN(n1713) );
  LVT_OAI21HSV2 U2177 ( .A1(n1715), .A2(n1714), .B(n1713), .ZN(n1188) );
  LVT_CLKNHSV2 U2189 ( .I(n577), .ZN(n1737) );
  LVT_OAI31HSV2 U2190 ( .A1(n1740), .A2(n2391), .A3(n1819), .B(n1738), .ZN(
        n1741) );
  LVT_INAND2HSV2 U2191 ( .A1(n3072), .B1(n1741), .ZN(n1744) );
  LVT_CLKNHSV2 U2192 ( .I(n1741), .ZN(n1742) );
  LVT_OAI21HSV2 U2193 ( .A1(n414), .A2(n1742), .B(C2_stall), .ZN(n1743) );
  LVT_OAI31HSV2 U2194 ( .A1(n1744), .A2(n1849), .A3(n1840), .B(n1743), .ZN(
        n1021) );
  LVT_INAND2HSV2 U2223 ( .A1(n3083), .B1(C1_N80), .ZN(n724) );
  LVT_CLKNHSV2 U2239 ( .I(n575), .ZN(n150) );
  LVT_INAND2HSV2 U2250 ( .A1(n1840), .B1(msg_C2_C1), .ZN(n1842) );
  LVT_OR4HSV0 U2251 ( .A1(n1898), .A2(n1842), .A3(n500), .A4(n2389), .Z(n1843)
         );
  LVT_OR4HSV0 U2252 ( .A1(n501), .A2(n2394), .A3(n1844), .A4(n1843), .Z(n496)
         );
  LVT_DQHSV2 C1_state_reg_2_ ( .D(n1127), .CK(clk), .Q(debugStateC1[2]) );
  LVT_EDGRNHSV1 C1_addr_reg_13_ ( .RN(C1_N80), .D(addr_C1_M[13]), .E(n3030), 
        .CK(clk), .Q(n1280), .QN(n1281) );
  LVT_EDGRNQHSV1 C1_addr_reg_4_ ( .RN(C1_N80), .D(addr_C1_M[4]), .E(n3030), 
        .CK(clk), .Q(C1_addr_4_) );
  LVT_EDGRNQHSV1 C1_addr_reg_15_ ( .RN(C1_N80), .D(addr_C1_M[15]), .E(n3031), 
        .CK(clk), .Q(C1_addr_15_) );
  LVT_DQHSV1 C1_state_reg_0_ ( .D(n1125), .CK(clk), .Q(debugStateC1[0]) );
  LVT_DQHSV1 C2_state_reg_2_ ( .D(n1077), .CK(clk), .Q(debugStateC2[2]) );
  LVT_DQHSV1 P2_addrToMem_reg_0_ ( .D(n1093), .CK(clk), .Q(addr_P2_C2[0]) );
  LVT_DQHSV1 C2_state_reg_1_ ( .D(n1076), .CK(clk), .Q(debugStateC2[1]) );
  LVT_DQHSV1 C2_state_reg_0_ ( .D(n1075), .CK(clk), .Q(debugStateC2[0]) );
  LVT_DHSV1 P2_addrToMem_reg_3_ ( .D(n1090), .CK(clk), .Q(n1290), .QN(n1916)
         );
  LVT_DQHSV1 mb_memEnB_reg ( .D(n1173), .CK(clk), .Q(en_M_C2) );
  LVT_DQHSV1 mb_memEnA_reg ( .D(n1210), .CK(clk), .Q(en_M_C1) );
  LVT_DQHSV1 P2_addrToMem_reg_14_ ( .D(n1079), .CK(clk), .Q(addr_P2_C2[14]) );
  LVT_DQHSV1 P2_addrToMem_reg_8_ ( .D(n1085), .CK(clk), .Q(addr_P2_C2[8]) );
  LVT_DQHSV1 P2_addrToMem_reg_7_ ( .D(n1086), .CK(clk), .Q(addr_P2_C2[7]) );
  LVT_DQHSV1 P2_addrToMem_reg_10_ ( .D(n1083), .CK(clk), .Q(addr_P2_C2[10]) );
  LVT_DQHSV1 P2_addrToMem_reg_4_ ( .D(n1089), .CK(clk), .Q(addr_P2_C2[4]) );
  LVT_DQHSV1 P2_addrToMem_reg_13_ ( .D(n1080), .CK(clk), .Q(addr_P2_C2[13]) );
  LVT_DQHSV1 P1_addrToMem_reg_15_ ( .D(n1128), .CK(clk), .Q(addr_P1_C1[15]) );
  LVT_DQHSV1 P1_addrToMem_reg_12_ ( .D(n1131), .CK(clk), .Q(addr_P1_C1[12]) );
  LVT_DQHSV1 P1_addrToMem_reg_13_ ( .D(n1130), .CK(clk), .Q(addr_P1_C1[13]) );
  LVT_DQHSV1 P1_addrToMem_reg_11_ ( .D(n1132), .CK(clk), .Q(addr_P1_C1[11]) );
  LVT_DQHSV1 P1_addrToMem_reg_3_ ( .D(n1140), .CK(clk), .Q(addr_P1_C1[3]) );
  LVT_EDGRNQHSV2 C2_addr_reg_10_ ( .RN(C1_N80), .D(addr_C2_M[10]), .E(n3028), 
        .CK(clk), .Q(C2_addr_10_) );
  LVT_EDGRNQHSV2 C2_addr_reg_0_ ( .RN(C1_N80), .D(addr_C2_M[0]), .E(n3028), 
        .CK(clk), .Q(C2_addr_0_) );
  LVT_EDGRNQHSV2 C2_addr_reg_8_ ( .RN(C1_N80), .D(addr_C2_M[8]), .E(n3028), 
        .CK(clk), .Q(C2_addr_8_) );
  LVT_EDGRNQHSV2 C2_addr_reg_2_ ( .RN(C1_N80), .D(addr_C2_M[2]), .E(n3028), 
        .CK(clk), .Q(C2_addr_2_) );
  LVT_EDGRNQHSV2 C2_addr_reg_4_ ( .RN(C1_N80), .D(addr_C2_M[4]), .E(n3028), 
        .CK(clk), .Q(C2_addr_4_) );
  LVT_EDGRNQHSV2 C2_addr_reg_11_ ( .RN(C1_N80), .D(addr_C2_M[11]), .E(n3029), 
        .CK(clk), .Q(C2_addr_11_) );
  LVT_EDGRNQHSV2 C2_addr_reg_14_ ( .RN(C1_N80), .D(addr_C2_M[14]), .E(n3028), 
        .CK(clk), .Q(C2_addr_14_) );
  LVT_EDGRNQHSV2 C2_addr_reg_7_ ( .RN(C1_N80), .D(addr_C2_M[7]), .E(n3029), 
        .CK(clk), .Q(C2_addr_7_) );
  LVT_EDGRNQHSV1 C1_addr_reg_9_ ( .RN(C1_N80), .D(addr_C1_M[9]), .E(n3030), 
        .CK(clk), .Q(C1_addr_9_) );
  LVT_EDGRNQHSV1 C1_addr_reg_10_ ( .RN(C1_N80), .D(addr_C1_M[10]), .E(n3031), 
        .CK(clk), .Q(C1_addr_10_) );
  LVT_EDGRNHSV1 C1_addr_reg_11_ ( .RN(C1_N80), .D(addr_C1_M[11]), .E(n3031), 
        .CK(clk), .Q(n1278), .QN(n1279) );
  LVT_EDGRNHSV1 C2_addr_reg_3_ ( .RN(C1_N80), .D(addr_C2_M[3]), .E(n3028), 
        .CK(clk), .Q(n1276), .QN(n1277) );
  LVT_EDGRNHSV1 C2_addr_reg_1_ ( .RN(C1_N80), .D(addr_C2_M[1]), .E(n3029), 
        .CK(clk), .Q(n1284), .QN(n1285) );
  LVT_EDGRNQHSV1 C2_addr_reg_15_ ( .RN(C1_N80), .D(addr_C2_M[15]), .E(n3028), 
        .CK(clk), .Q(C2_addr_15_) );
  LVT_EDGRNQHSV1 C2_addr_reg_12_ ( .RN(C1_N80), .D(addr_C2_M[12]), .E(n3029), 
        .CK(clk), .Q(C2_addr_12_) );
  LVT_EDGRNQHSV1 C2_addr_reg_9_ ( .RN(C1_N80), .D(addr_C2_M[9]), .E(n3029), 
        .CK(clk), .Q(C2_addr_9_) );
  LVT_EDGRNQHSV1 C2_addr_reg_6_ ( .RN(C1_N80), .D(addr_C2_M[6]), .E(n3029), 
        .CK(clk), .Q(C2_addr_6_) );
  LVT_EDGRNQHSV1 C2_addr_reg_13_ ( .RN(C1_N80), .D(addr_C2_M[13]), .E(n3029), 
        .CK(clk), .Q(C2_addr_13_) );
  LVT_EDGRNQHSV1 C2_addr_reg_5_ ( .RN(C1_N80), .D(addr_C2_M[5]), .E(n3029), 
        .CK(clk), .Q(C2_addr_5_) );
  LVT_DQHSV1 P2_addrToMem_reg_12_ ( .D(n1081), .CK(clk), .Q(addr_P2_C2[12]) );
  LVT_DQHSV1 P1_addrToMem_reg_4_ ( .D(n1139), .CK(clk), .Q(addr_P1_C1[4]) );
  LVT_DQHSV1 C2_state_reg_3_ ( .D(n1190), .CK(clk), .Q(debugStateC2[3]) );
  LVT_DQHSV1 C1_state_reg_3_ ( .D(n1209), .CK(clk), .Q(debugStateC1[3]) );
  LVT_DQHSV1 C1_state_reg_1_ ( .D(n1126), .CK(clk), .Q(debugStateC1[1]) );
  LVT_OAI211HSV1 U2040 ( .A1(n2997), .A2(n2954), .B(n3017), .C(n2953), .ZN(
        n725) );
  CLKNHSV0 U2043 ( .I(addr_C1_M[8]), .ZN(n2593) );
  CLKNHSV0 U2044 ( .I(addr_C1_M[13]), .ZN(n2594) );
  HVT_OAI22HSV0 U2047 ( .A1(n2593), .A2(addr_P1_C1[8]), .B1(n2594), .B2(
        addr_P1_C1[13]), .ZN(n2595) );
  AOI221HSV0 U2048 ( .A1(n2593), .A2(addr_P1_C1[8]), .B1(addr_P1_C1[13]), .B2(
        n2594), .C(n2595), .ZN(n2674) );
  LVT_OR2HSV1 U2051 ( .A1(n2834), .A2(n2686), .Z(n2932) );
  AND2HSV0 U2052 ( .A1(n2840), .A2(n2955), .Z(n2596) );
  AOI21HSV0 U2055 ( .A1(n2862), .A2(n2853), .B(en_M_C2), .ZN(n2597) );
  AOI211HSV0 U2057 ( .A1(n2849), .A2(n2596), .B(n3071), .C(n2597), .ZN(n737)
         );
  HVT_INOR2HSV0 U2058 ( .A1(C2_stall), .B1(n534), .ZN(n3069) );
  LVT_INHSV2 U2059 ( .I(addr_C2_C1[3]), .ZN(n2598) );
  LVT_INHSV2 U2068 ( .I(addr_C2_C1[7]), .ZN(n2599) );
  LVT_AOI22HSV2 U2069 ( .A1(C1_addr_3_), .A2(n2598), .B1(C1_addr_7_), .B2(
        n2599), .ZN(n2600) );
  LVT_OAI221HSV1 U2070 ( .A1(n2598), .A2(C1_addr_3_), .B1(n2599), .B2(
        C1_addr_7_), .C(n2600), .ZN(n2634) );
  CLKNHSV0 U2071 ( .I(addr_C1_M[12]), .ZN(n2601) );
  CLKNHSV0 U2072 ( .I(addr_C1_M[11]), .ZN(n2602) );
  HVT_OAI22HSV0 U2074 ( .A1(n2601), .A2(addr_P1_C1[12]), .B1(n2602), .B2(
        addr_P1_C1[11]), .ZN(n2603) );
  AOI221HSV0 U2077 ( .A1(n2601), .A2(addr_P1_C1[12]), .B1(addr_P1_C1[11]), 
        .B2(n2602), .C(n2603), .ZN(n2675) );
  HVT_NAND3HSV0 U2078 ( .A1(n2929), .A2(en_M_C1), .A3(n3049), .ZN(n2965) );
  HVT_INAND3HSV0 U2085 ( .A1(C1_stall), .B1(n3044), .B2(n1555), .ZN(n2970) );
  HVT_OR2HSV0 U2088 ( .A1(debugStateC1[2]), .A2(debugStateC1[3]), .Z(n2930) );
  HVT_INAND2HSV0 U2090 ( .A1(n3071), .B1(n2956), .ZN(n1844) );
  LVT_INOR3HSV2 U2091 ( .A1(n2773), .B1(debugStateC2[1]), .B2(n2783), .ZN(
        n3070) );
  HVT_OR4HSV0 U2092 ( .A1(n1898), .A2(n2861), .A3(n3083), .A4(n500), .Z(n2809)
         );
  LVT_NOR4HSV2 U2093 ( .A1(n2681), .A2(n2680), .A3(n2679), .A4(n2678), .ZN(
        n2604) );
  HVT_NAND3HSV0 U2095 ( .A1(n2604), .A2(n2676), .A3(n2677), .ZN(n2605) );
  LVT_NOR4HSV2 U2096 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(
        n2606) );
  HVT_NAND3HSV0 U2097 ( .A1(n2606), .A2(n2674), .A3(n2675), .ZN(n2607) );
  LVT_OAI21HSV2 U2103 ( .A1(n2605), .A2(n2607), .B(n1789), .ZN(n2737) );
  HVT_INOR2HSV0 U2105 ( .A1(n2926), .B1(n2927), .ZN(n3041) );
  HVT_IOA21HSV0 U2106 ( .A1(en_M_C1), .A2(n3045), .B(n600), .ZN(n2512) );
  HVT_OAI211HSV0 U2107 ( .A1(n3023), .A2(n3072), .B(n3070), .C(n3022), .ZN(
        n2608) );
  HVT_INAND3HSV0 U2108 ( .A1(n3037), .B1(n3024), .B2(n2608), .ZN(n2609) );
  HVT_NAND3HSV0 U2110 ( .A1(n3026), .A2(n3025), .A3(n513), .ZN(n2610) );
  AOI211HSV0 U2111 ( .A1(n3074), .A2(n3069), .B(n2609), .C(n2610), .ZN(n3033)
         );
  LVT_INAND3HSV2 U2112 ( .A1(n2863), .B1(n3100), .B2(n3078), .ZN(n3003) );
  HVT_INAND3HSV0 U2113 ( .A1(n2931), .B1(n2834), .B2(n3064), .ZN(n2611) );
  HVT_OAI211HSV0 U2114 ( .A1(n2929), .A2(n1672), .B(n2964), .C(n2611), .ZN(
        n2612) );
  HVT_NOR2HSV0 U2118 ( .A1(n2968), .A2(n2612), .ZN(n631) );
  CLKNHSV0 U2120 ( .I(en_M_C2), .ZN(n2613) );
  CLKNHSV0 U2121 ( .I(n1898), .ZN(n2614) );
  AOI21HSV0 U2122 ( .A1(n2854), .A2(n2614), .B(n3004), .ZN(n2615) );
  HVT_INOR2HSV0 U2123 ( .A1(n522), .B1(n2853), .ZN(n2616) );
  AOI211HSV0 U2124 ( .A1(n3084), .A2(n2613), .B(n2615), .C(n2616), .ZN(n511)
         );
  HVT_INAND3HSV0 U2125 ( .A1(n465), .B1(n2987), .B2(n3061), .ZN(n1789) );
  CLKNHSV0 U2126 ( .I(addr_C1_M[14]), .ZN(n2617) );
  CLKNHSV0 U2127 ( .I(addr_C1_M[7]), .ZN(n2618) );
  HVT_OAI22HSV0 U2128 ( .A1(n2617), .A2(addr_P1_C1[14]), .B1(n2618), .B2(
        addr_P1_C1[7]), .ZN(n2619) );
  AOI221HSV0 U2129 ( .A1(n2617), .A2(addr_P1_C1[14]), .B1(addr_P1_C1[7]), .B2(
        n2618), .C(n2619), .ZN(n2676) );
  AO32HSV0 U2130 ( .A1(n2928), .A2(n3061), .A3(n2932), .B1(n2928), .B2(en_M_C1), .Z(n2620) );
  HVT_NAND4HSV0 U2131 ( .A1(n2966), .A2(n2970), .A3(n2858), .A4(n2620), .ZN(
        n1568) );
  HVT_INAND2HSV0 U2132 ( .A1(n2852), .B1(en_M_C2), .ZN(n522) );
  CLKNAND2HSV0 U2133 ( .A1(n2952), .A2(n431), .ZN(n2621) );
  HVT_NOR3HSV0 U2134 ( .A1(n3009), .A2(n3046), .A3(n2621), .ZN(n1811) );
  HVT_OR2HSV0 U2135 ( .A1(n2859), .A2(n2930), .Z(n600) );
  HVT_INOR3HSV0 U2140 ( .A1(debugStateC2[0]), .B1(debugStateC2[1]), .B2(n2938), 
        .ZN(n3037) );
  LVT_XNOR2HSV1 U2141 ( .A1(addr_C2_C1[15]), .A2(C1_addr_15_), .ZN(n2625) );
  LVT_XNOR2HSV1 U2146 ( .A1(addr_C2_C1[2]), .A2(C1_addr_2_), .ZN(n2624) );
  LVT_XNOR2HSV1 U2151 ( .A1(addr_C2_C1[5]), .A2(C1_addr_5_), .ZN(n2623) );
  LVT_XNOR2HSV1 U2156 ( .A1(addr_C2_C1[1]), .A2(C1_addr_1_), .ZN(n2622) );
  LVT_NAND4HSV2 U2159 ( .A1(n2625), .A2(n2624), .A3(n2623), .A4(n2622), .ZN(
        n2631) );
  LVT_XNOR2HSV1 U2165 ( .A1(addr_C2_C1[14]), .A2(C1_addr_14_), .ZN(n2629) );
  LVT_XNOR2HSV1 U2166 ( .A1(addr_C2_C1[0]), .A2(C1_addr_0_), .ZN(n2628) );
  LVT_XNOR2HSV1 U2167 ( .A1(addr_C2_C1[11]), .A2(n1278), .ZN(n2627) );
  LVT_XNOR2HSV1 U2170 ( .A1(addr_C2_C1[9]), .A2(C1_addr_9_), .ZN(n2626) );
  LVT_NAND4HSV2 U2175 ( .A1(n2629), .A2(n2628), .A3(n2627), .A4(n2626), .ZN(
        n2630) );
  LVT_NOR2HSV2 U2178 ( .A1(n2631), .A2(n2630), .ZN(n2642) );
  LVT_XOR2HSV0 U2179 ( .A1(addr_C2_C1[4]), .A2(C1_addr_4_), .Z(n2633) );
  LVT_XOR2HSV0 U2180 ( .A1(addr_C2_C1[8]), .A2(C1_addr_8_), .Z(n2632) );
  LVT_NOR3HSV2 U2181 ( .A1(n2634), .A2(n2633), .A3(n2632), .ZN(n2641) );
  LVT_XNOR2HSV1 U2182 ( .A1(n1296), .A2(addr_C2_C1[12]), .ZN(n2636) );
  LVT_XNOR2HSV1 U2183 ( .A1(C1_addr_10_), .A2(n1293), .ZN(n2635) );
  LVT_NAND3HSV2 U2184 ( .A1(n2636), .A2(msg_C2_C1), .A3(n2635), .ZN(n2639) );
  LVT_XOR2HSV0 U2185 ( .A1(n1280), .A2(addr_C2_C1[13]), .Z(n2638) );
  LVT_XOR2HSV0 U2186 ( .A1(addr_C2_C1[6]), .A2(C1_addr_6_), .Z(n2637) );
  LVT_NOR3HSV2 U2187 ( .A1(n2639), .A2(n2638), .A3(n2637), .ZN(n2640) );
  LVT_NAND3HSV2 U2188 ( .A1(n2642), .A2(n2641), .A3(n2640), .ZN(n2643) );
  LVT_INHSV2 U2195 ( .I(rm_C2_C1), .ZN(n2843) );
  LVT_NOR2HSV2 U2196 ( .A1(n2643), .A2(n2843), .ZN(n2969) );
  LVT_INHSV2 U2197 ( .I(wm_C2_C1), .ZN(n2483) );
  LVT_NOR2HSV2 U2198 ( .A1(n2643), .A2(n2483), .ZN(n2864) );
  LVT_NOR2HSV4 U2199 ( .A1(n2969), .A2(n2864), .ZN(n2959) );
  LVT_INOR2HSV1 U2200 ( .A1(rw_P1_C1[1]), .B1(rw_P1_C1[0]), .ZN(n3065) );
  LVT_NAND2HSV2 U2201 ( .A1(n2959), .A2(n3065), .ZN(n592) );
  LVT_INHSV2 U2202 ( .I(debugStateC1[1]), .ZN(n2855) );
  LVT_NAND2HSV2 U2203 ( .A1(n2855), .A2(debugStateC1[0]), .ZN(n2927) );
  LVT_NOR2HSV2 U2204 ( .A1(n2930), .A2(n2927), .ZN(n3068) );
  LVT_INHSV2 U2205 ( .I(n3068), .ZN(n2865) );
  LVT_NOR2HSV2 U2206 ( .A1(n592), .A2(n2865), .ZN(n3056) );
  LVT_XOR2HSV0 U2207 ( .A1(C1_addr_8_), .A2(addr_P1_C1[8]), .Z(n2645) );
  LVT_XOR2HSV0 U2208 ( .A1(C1_addr_7_), .A2(addr_P1_C1[7]), .Z(n2644) );
  LVT_NOR2HSV2 U2209 ( .A1(n2645), .A2(n2644), .ZN(n2655) );
  LVT_XOR2HSV0 U2210 ( .A1(C1_addr_2_), .A2(addr_P1_C1[2]), .Z(n2647) );
  LVT_XOR2HSV0 U2211 ( .A1(C1_addr_6_), .A2(addr_P1_C1[6]), .Z(n2646) );
  LVT_NOR2HSV2 U2212 ( .A1(n2647), .A2(n2646), .ZN(n2654) );
  LVT_XOR2HSV0 U2213 ( .A1(addr_P1_C1[9]), .A2(C1_addr_9_), .Z(n2649) );
  LVT_XOR2HSV0 U2214 ( .A1(addr_P1_C1[10]), .A2(C1_addr_10_), .Z(n2648) );
  LVT_NOR2HSV2 U2215 ( .A1(n2649), .A2(n2648), .ZN(n2653) );
  LVT_XOR2HSV0 U2216 ( .A1(C1_addr_14_), .A2(addr_P1_C1[14]), .Z(n2651) );
  LVT_XOR2HSV0 U2217 ( .A1(n1278), .A2(addr_P1_C1[11]), .Z(n2650) );
  LVT_NOR2HSV2 U2218 ( .A1(n2651), .A2(n2650), .ZN(n2652) );
  LVT_NAND4HSV2 U2219 ( .A1(n2655), .A2(n2654), .A3(n2653), .A4(n2652), .ZN(
        n2669) );
  LVT_XOR2HSV0 U2220 ( .A1(C1_addr_5_), .A2(addr_P1_C1[5]), .Z(n2657) );
  LVT_XOR2HSV0 U2221 ( .A1(C1_addr_1_), .A2(addr_P1_C1[1]), .Z(n2656) );
  LVT_NOR2HSV2 U2222 ( .A1(n2657), .A2(n2656), .ZN(n2667) );
  LVT_XOR2HSV0 U2224 ( .A1(n1280), .A2(addr_P1_C1[13]), .Z(n2659) );
  LVT_XOR2HSV0 U2225 ( .A1(n1296), .A2(addr_P1_C1[12]), .Z(n2658) );
  LVT_NOR2HSV2 U2226 ( .A1(n2659), .A2(n2658), .ZN(n2666) );
  LVT_XOR2HSV0 U2227 ( .A1(C1_addr_3_), .A2(addr_P1_C1[3]), .Z(n2661) );
  LVT_XOR2HSV0 U2228 ( .A1(C1_addr_4_), .A2(addr_P1_C1[4]), .Z(n2660) );
  LVT_NOR2HSV2 U2229 ( .A1(n2661), .A2(n2660), .ZN(n2665) );
  LVT_XOR2HSV0 U2230 ( .A1(C1_addr_0_), .A2(addr_P1_C1[0]), .Z(n2663) );
  LVT_XOR2HSV0 U2231 ( .A1(C1_addr_15_), .A2(addr_P1_C1[15]), .Z(n2662) );
  LVT_NOR2HSV2 U2232 ( .A1(n2663), .A2(n2662), .ZN(n2664) );
  LVT_NAND4HSV2 U2233 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(
        n2668) );
  LVT_NOR2HSV2 U2234 ( .A1(n2669), .A2(n2668), .ZN(n2958) );
  LVT_INAND2HSV2 U2235 ( .A1(debugStateC1[2]), .B1(debugStateC1[3]), .ZN(n2671) );
  LVT_CLKNAND2HSV1 U2236 ( .A1(debugStateC1[0]), .A2(debugStateC1[1]), .ZN(
        n2859) );
  LVT_NOR2HSV2 U2237 ( .A1(n2671), .A2(n2859), .ZN(n3054) );
  LVT_INHSV2 U2238 ( .I(n3054), .ZN(n2957) );
  LVT_AOI21HSV2 U2240 ( .A1(n2958), .A2(n2957), .B(rw_P1_C1[1]), .ZN(n3053) );
  LVT_NAND2HSV2 U2241 ( .A1(n2959), .A2(n3053), .ZN(n2963) );
  LVT_INAND2HSV2 U2242 ( .A1(debugStateC1[0]), .B1(n2855), .ZN(n2686) );
  LVT_NOR2HSV2 U2243 ( .A1(n2686), .A2(n2671), .ZN(n3055) );
  LVT_INHSV2 U2244 ( .I(n3055), .ZN(n591) );
  LVT_OAI22HSV2 U2245 ( .A1(n2963), .A2(n591), .B1(rw_P1_C1[1]), .B2(n2957), 
        .ZN(n2011) );
  LVT_INHSV2 U2246 ( .I(n2963), .ZN(n2670) );
  LVT_NAND2HSV0 U2247 ( .A1(n2670), .A2(n3068), .ZN(n2858) );
  LVT_INAND2HSV2 U2248 ( .A1(debugStateC1[0]), .B1(debugStateC1[1]), .ZN(n2931) );
  LVT_NOR2HSV2 U2249 ( .A1(n2931), .A2(n2671), .ZN(n2743) );
  LVT_NOR2HSV2 U2253 ( .A1(n2927), .A2(n2671), .ZN(n3060) );
  LVT_XOR2HSV0 U2254 ( .A1(addr_C1_M[10]), .A2(addr_P1_C1[10]), .Z(n2673) );
  LVT_XOR2HSV0 U2255 ( .A1(addr_C1_M[9]), .A2(addr_P1_C1[9]), .Z(n2672) );
  LVT_NOR2HSV2 U2256 ( .A1(n2673), .A2(n2672), .ZN(n2677) );
  LVT_XOR2HSV0 U2257 ( .A1(addr_C1_M[0]), .A2(addr_P1_C1[0]), .Z(n2679) );
  LVT_XOR2HSV0 U2258 ( .A1(addr_C1_M[15]), .A2(addr_P1_C1[15]), .Z(n2678) );
  LVT_XOR2HSV0 U2259 ( .A1(addr_C1_M[5]), .A2(addr_P1_C1[5]), .Z(n2681) );
  LVT_XOR2HSV0 U2260 ( .A1(addr_C1_M[6]), .A2(addr_P1_C1[6]), .Z(n2680) );
  LVT_XOR2HSV0 U2261 ( .A1(addr_C1_M[2]), .A2(addr_P1_C1[2]), .Z(n2683) );
  LVT_XOR2HSV0 U2262 ( .A1(addr_C1_M[3]), .A2(addr_P1_C1[3]), .Z(n2682) );
  LVT_XOR2HSV0 U2263 ( .A1(addr_C1_M[1]), .A2(addr_P1_C1[1]), .Z(n2685) );
  LVT_XOR2HSV0 U2264 ( .A1(addr_C1_M[4]), .A2(addr_P1_C1[4]), .Z(n2684) );
  LVT_INOR2HSV1 U2265 ( .A1(debugStateC1[2]), .B1(debugStateC1[3]), .ZN(n2926)
         );
  LVT_INOR2HSV1 U2266 ( .A1(n2926), .B1(n2931), .ZN(n2740) );
  LVT_CLKNAND2HSV0 U2267 ( .A1(debugStateC1[3]), .A2(debugStateC1[2]), .ZN(
        n2834) );
  LVT_NOR2HSV2 U2268 ( .A1(n2927), .A2(n2834), .ZN(n2835) );
  LVT_NOR2HSV2 U2269 ( .A1(n2740), .A2(n2835), .ZN(n3063) );
  LVT_INAND2HSV2 U2270 ( .A1(n2859), .B1(n2926), .ZN(n639) );
  LVT_CLKAND2HSV2 U2271 ( .A1(n3063), .A2(n639), .Z(n3061) );
  LVT_INAND2HSV2 U2272 ( .A1(n3060), .B1(n2932), .ZN(n465) );
  LVT_INHSV2 U2273 ( .I(n2743), .ZN(n2987) );
  LVT_NAND2HSV2 U2274 ( .A1(n2737), .A2(en_M_C1), .ZN(n1674) );
  LVT_OAI21HSV0 U2275 ( .A1(n2743), .A2(n3060), .B(n1674), .ZN(n2687) );
  LVT_NAND3HSV0 U2276 ( .A1(n2858), .A2(n2687), .A3(n2932), .ZN(n2688) );
  LVT_AOI211HSV0 U2277 ( .A1(msg_C1_C2), .A2(n3056), .B(n2011), .C(n2688), 
        .ZN(n1657) );
  LVT_XNOR2HSV1 U2278 ( .A1(addr_C1_C2[14]), .A2(C2_addr_14_), .ZN(n2692) );
  LVT_XNOR2HSV1 U2279 ( .A1(addr_C1_C2[7]), .A2(C2_addr_7_), .ZN(n2691) );
  LVT_XNOR2HSV1 U2280 ( .A1(addr_C1_C2[10]), .A2(C2_addr_10_), .ZN(n2690) );
  LVT_XNOR2HSV1 U2281 ( .A1(C2_addr_6_), .A2(addr_C1_C2[6]), .ZN(n2689) );
  LVT_NAND4HSV2 U2282 ( .A1(n2692), .A2(n2691), .A3(n2690), .A4(n2689), .ZN(
        n2698) );
  LVT_XNOR2HSV1 U2283 ( .A1(addr_C1_C2[8]), .A2(C2_addr_8_), .ZN(n2696) );
  LVT_XNOR2HSV1 U2284 ( .A1(addr_C1_C2[11]), .A2(C2_addr_11_), .ZN(n2695) );
  LVT_XNOR2HSV1 U2285 ( .A1(addr_C1_C2[0]), .A2(C2_addr_0_), .ZN(n2694) );
  LVT_XNOR2HSV1 U2286 ( .A1(addr_C1_C2[9]), .A2(C2_addr_9_), .ZN(n2693) );
  LVT_NAND4HSV2 U2287 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(
        n2697) );
  LVT_NOR2HSV2 U2288 ( .A1(n2698), .A2(n2697), .ZN(n2711) );
  LVT_XNOR2HSV1 U2289 ( .A1(n1276), .A2(addr_C1_C2[3]), .ZN(n2700) );
  LVT_XNOR2HSV1 U2290 ( .A1(addr_C1_C2[15]), .A2(C2_addr_15_), .ZN(n2699) );
  LVT_NAND3HSV2 U2291 ( .A1(n2700), .A2(msg_C1_C2), .A3(n2699), .ZN(n2703) );
  LVT_XOR2HSV0 U2292 ( .A1(n1284), .A2(addr_C1_C2[1]), .Z(n2702) );
  LVT_XOR2HSV0 U2293 ( .A1(addr_C1_C2[13]), .A2(C2_addr_13_), .Z(n2701) );
  LVT_NOR3HSV2 U2294 ( .A1(n2703), .A2(n2702), .A3(n2701), .ZN(n2710) );
  LVT_XNOR2HSV1 U2295 ( .A1(addr_C1_C2[2]), .A2(C2_addr_2_), .ZN(n2705) );
  LVT_XNOR2HSV1 U2296 ( .A1(addr_C1_C2[12]), .A2(C2_addr_12_), .ZN(n2704) );
  LVT_NAND2HSV2 U2297 ( .A1(n2705), .A2(n2704), .ZN(n2708) );
  LVT_XOR2HSV0 U2298 ( .A1(addr_C1_C2[5]), .A2(C2_addr_5_), .Z(n2707) );
  LVT_XOR2HSV0 U2299 ( .A1(addr_C1_C2[4]), .A2(C2_addr_4_), .Z(n2706) );
  LVT_NOR3HSV2 U2300 ( .A1(n2708), .A2(n2707), .A3(n2706), .ZN(n2709) );
  LVT_NAND3HSV2 U2301 ( .A1(n2711), .A2(n2710), .A3(n2709), .ZN(n2713) );
  LVT_INHSV2 U2302 ( .I(wm_C1_C2), .ZN(n2712) );
  LVT_NOR2HSV2 U2303 ( .A1(n2713), .A2(n2712), .ZN(n3023) );
  LVT_INHSV2 U2304 ( .I(rm_C1_C2), .ZN(n2780) );
  LVT_NOR2HSV2 U2305 ( .A1(n2713), .A2(n2780), .ZN(n3018) );
  LVT_NOR2HSV4 U2306 ( .A1(n3023), .A2(n3018), .ZN(n3078) );
  LVT_NAND2HSV2 U2307 ( .A1(n3078), .A2(rw_P2_C2[0]), .ZN(n2849) );
  LVT_INHSV2 U2308 ( .I(rw_P2_C2[1]), .ZN(n3100) );
  LVT_INAND2HSV2 U2309 ( .A1(debugStateC2[2]), .B1(debugStateC2[0]), .ZN(n2783) );
  LVT_INHSV2 U2310 ( .I(debugStateC2[3]), .ZN(n2773) );
  LVT_OAI21HSV2 U2311 ( .A1(n2849), .A2(n3100), .B(n3070), .ZN(n431) );
  LVT_INHSV2 U2312 ( .I(rw_P1_C1[0]), .ZN(n3066) );
  LVT_AND2HSV2 U2313 ( .A1(n3053), .A2(n3066), .Z(n3043) );
  LVT_NAND3HSV2 U2314 ( .A1(n3043), .A2(n2959), .A3(n3055), .ZN(n2778) );
  LVT_INHSV2 U2315 ( .I(n2778), .ZN(n3042) );
  LVT_XNOR2HSV0 U2316 ( .A1(allowReadAddr_C2_C1[10]), .A2(addr_P1_C1[10]), 
        .ZN(n2717) );
  LVT_XNOR2HSV0 U2317 ( .A1(allowReadAddr_C2_C1[6]), .A2(addr_P1_C1[6]), .ZN(
        n2716) );
  LVT_XNOR2HSV0 U2318 ( .A1(allowReadAddr_C2_C1[2]), .A2(addr_P1_C1[2]), .ZN(
        n2715) );
  LVT_XNOR2HSV0 U2319 ( .A1(allowReadAddr_C2_C1[9]), .A2(addr_P1_C1[9]), .ZN(
        n2714) );
  LVT_NAND4HSV2 U2320 ( .A1(n2717), .A2(n2716), .A3(n2715), .A4(n2714), .ZN(
        n2723) );
  LVT_XNOR2HSV0 U2321 ( .A1(allowReadAddr_C2_C1[7]), .A2(addr_P1_C1[7]), .ZN(
        n2721) );
  LVT_XNOR2HSV0 U2322 ( .A1(allowReadAddr_C2_C1[11]), .A2(addr_P1_C1[11]), 
        .ZN(n2720) );
  LVT_XNOR2HSV0 U2323 ( .A1(allowReadAddr_C2_C1[4]), .A2(addr_P1_C1[4]), .ZN(
        n2719) );
  LVT_XNOR2HSV0 U2324 ( .A1(allowReadAddr_C2_C1[3]), .A2(addr_P1_C1[3]), .ZN(
        n2718) );
  LVT_NAND4HSV2 U2325 ( .A1(n2721), .A2(n2720), .A3(n2719), .A4(n2718), .ZN(
        n2722) );
  LVT_NOR2HSV2 U2326 ( .A1(n2723), .A2(n2722), .ZN(n2736) );
  LVT_XNOR2HSV0 U2327 ( .A1(allowReadAddr_C2_C1[5]), .A2(addr_P1_C1[5]), .ZN(
        n2727) );
  LVT_XNOR2HSV0 U2328 ( .A1(allowReadAddr_C2_C1[1]), .A2(addr_P1_C1[1]), .ZN(
        n2726) );
  LVT_XNOR2HSV0 U2329 ( .A1(allowReadAddr_C2_C1[0]), .A2(addr_P1_C1[0]), .ZN(
        n2725) );
  LVT_XNOR2HSV0 U2330 ( .A1(allowReadAddr_C2_C1[12]), .A2(addr_P1_C1[12]), 
        .ZN(n2724) );
  LVT_AND4HSV1 U2331 ( .A1(n2727), .A2(n2726), .A3(n2725), .A4(n2724), .Z(
        n2735) );
  LVT_XNOR2HSV0 U2332 ( .A1(allowReadAddr_C2_C1[14]), .A2(addr_P1_C1[14]), 
        .ZN(n2729) );
  LVT_XNOR2HSV0 U2333 ( .A1(allowReadAddr_C2_C1[8]), .A2(addr_P1_C1[8]), .ZN(
        n2728) );
  LVT_INHSV2 U2334 ( .I(allowRead_C2_C1), .ZN(n2810) );
  LVT_NAND3HSV2 U2335 ( .A1(n2729), .A2(n2728), .A3(n2810), .ZN(n2733) );
  LVT_XNOR2HSV0 U2336 ( .A1(allowReadAddr_C2_C1[15]), .A2(addr_P1_C1[15]), 
        .ZN(n2731) );
  LVT_XNOR2HSV0 U2337 ( .A1(allowReadAddr_C2_C1[13]), .A2(addr_P1_C1[13]), 
        .ZN(n2730) );
  LVT_CLKNAND2HSV1 U2338 ( .A1(n2731), .A2(n2730), .ZN(n2732) );
  LVT_NOR2HSV2 U2339 ( .A1(n2733), .A2(n2732), .ZN(n2734) );
  LVT_NAND3HSV2 U2340 ( .A1(n2736), .A2(n2735), .A3(n2734), .ZN(n2929) );
  LVT_NAND2HSV2 U2341 ( .A1(n3042), .A2(n2929), .ZN(n2971) );
  LVT_INAND2HSV0 U2342 ( .A1(n2737), .B1(en_M_C1), .ZN(n624) );
  LVT_CLKNHSV0 U2343 ( .I(n3060), .ZN(n2738) );
  LVT_CLKNHSV0 U2344 ( .I(rw_P1_C1[1]), .ZN(n3067) );
  LVT_NAND3HSV1 U2345 ( .A1(n3054), .A2(rw_P1_C1[0]), .A3(n3067), .ZN(n1672)
         );
  LVT_OAI21HSV0 U2346 ( .A1(n2738), .A2(en_M_C1), .B(n1672), .ZN(n2739) );
  LVT_AOI21HSV0 U2347 ( .A1(n624), .A2(n2835), .B(n2739), .ZN(n2742) );
  LVT_CLKNHSV0 U2348 ( .I(n1674), .ZN(n3058) );
  LVT_OAI21HSV0 U2349 ( .A1(n2743), .A2(n2740), .B(n3058), .ZN(n2741) );
  LVT_NAND3HSV0 U2350 ( .A1(n2971), .A2(n2742), .A3(n2741), .ZN(n1564) );
  LVT_NOR2HSV2 U2351 ( .A1(n2963), .A2(n3066), .ZN(n2745) );
  LVT_NAND2HSV2 U2352 ( .A1(n2745), .A2(n3055), .ZN(n2833) );
  LVT_INOR2HSV0 U2353 ( .A1(n2833), .B1(n2743), .ZN(n3052) );
  LVT_CLKNHSV0 U2354 ( .I(n3052), .ZN(n2744) );
  LVT_AOI211HSV0 U2355 ( .A1(n3068), .A2(n2745), .B(n3054), .C(n2744), .ZN(
        n1679) );
  LVT_INHSV2 U2356 ( .I(rw_P2_C2[0]), .ZN(n3076) );
  LVT_NAND2HSV2 U2357 ( .A1(rw_P2_C2[1]), .A2(n3076), .ZN(n2847) );
  LVT_INHSV2 U2358 ( .I(n2847), .ZN(n3072) );
  LVT_NAND2HSV2 U2359 ( .A1(n3078), .A2(n3072), .ZN(n694) );
  LVT_INHSV2 U2360 ( .I(n3070), .ZN(n444) );
  LVT_NOR2HSV2 U2361 ( .A1(n694), .A2(n444), .ZN(n3047) );
  LVT_CLKNHSV0 U2362 ( .I(n3047), .ZN(n420) );
  LVT_XOR2HSV0 U2363 ( .A1(C2_addr_11_), .A2(addr_P2_C2[11]), .Z(n2747) );
  LVT_XOR2HSV0 U2364 ( .A1(C2_addr_7_), .A2(addr_P2_C2[7]), .Z(n2746) );
  LVT_NOR2HSV2 U2365 ( .A1(n2747), .A2(n2746), .ZN(n2757) );
  LVT_XOR2HSV0 U2366 ( .A1(n1284), .A2(addr_P2_C2[1]), .Z(n2749) );
  LVT_XOR2HSV0 U2367 ( .A1(n1276), .A2(n1290), .Z(n2748) );
  LVT_NOR2HSV2 U2368 ( .A1(n2749), .A2(n2748), .ZN(n2756) );
  LVT_XOR2HSV0 U2369 ( .A1(C2_addr_13_), .A2(addr_P2_C2[13]), .Z(n2751) );
  LVT_XOR2HSV0 U2370 ( .A1(C2_addr_4_), .A2(addr_P2_C2[4]), .Z(n2750) );
  LVT_NOR2HSV2 U2371 ( .A1(n2751), .A2(n2750), .ZN(n2755) );
  LVT_XOR2HSV0 U2372 ( .A1(C2_addr_6_), .A2(addr_P2_C2[6]), .Z(n2753) );
  LVT_XOR2HSV0 U2373 ( .A1(C2_addr_0_), .A2(addr_P2_C2[0]), .Z(n2752) );
  LVT_NOR2HSV2 U2374 ( .A1(n2753), .A2(n2752), .ZN(n2754) );
  LVT_NAND4HSV2 U2375 ( .A1(n2757), .A2(n2756), .A3(n2755), .A4(n2754), .ZN(
        n2771) );
  LVT_XOR2HSV0 U2376 ( .A1(C2_addr_8_), .A2(addr_P2_C2[8]), .Z(n2759) );
  LVT_XOR2HSV0 U2377 ( .A1(C2_addr_14_), .A2(addr_P2_C2[14]), .Z(n2758) );
  LVT_NOR2HSV2 U2378 ( .A1(n2759), .A2(n2758), .ZN(n2769) );
  LVT_XOR2HSV0 U2379 ( .A1(C2_addr_2_), .A2(addr_P2_C2[2]), .Z(n2761) );
  LVT_XOR2HSV0 U2380 ( .A1(C2_addr_5_), .A2(addr_P2_C2[5]), .Z(n2760) );
  LVT_NOR2HSV2 U2381 ( .A1(n2761), .A2(n2760), .ZN(n2768) );
  LVT_XOR2HSV0 U2382 ( .A1(C2_addr_9_), .A2(addr_P2_C2[9]), .Z(n2763) );
  LVT_XOR2HSV0 U2383 ( .A1(C2_addr_10_), .A2(addr_P2_C2[10]), .Z(n2762) );
  LVT_NOR2HSV2 U2384 ( .A1(n2763), .A2(n2762), .ZN(n2767) );
  LVT_XOR2HSV0 U2385 ( .A1(C2_addr_15_), .A2(addr_P2_C2[15]), .Z(n2765) );
  LVT_XOR2HSV0 U2386 ( .A1(C2_addr_12_), .A2(addr_P2_C2[12]), .Z(n2764) );
  LVT_NOR2HSV2 U2387 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  LVT_NAND4HSV2 U2388 ( .A1(n2769), .A2(n2768), .A3(n2767), .A4(n2766), .ZN(
        n2770) );
  LVT_NOR2HSV2 U2389 ( .A1(n2771), .A2(n2770), .ZN(n2863) );
  LVT_AND2HSV2 U2390 ( .A1(n2863), .A2(n3100), .Z(n3077) );
  LVT_INHSV2 U2391 ( .I(n3077), .ZN(n2772) );
  LVT_CLKNAND2HSV2 U2392 ( .A1(n3078), .A2(n2772), .ZN(n2840) );
  LVT_NOR2HSV2 U2393 ( .A1(n2773), .A2(debugStateC2[2]), .ZN(n2774) );
  LVT_AND2HSV2 U2394 ( .A1(debugStateC2[0]), .A2(debugStateC2[1]), .Z(n2844)
         );
  LVT_NAND2HSV2 U2395 ( .A1(n2774), .A2(n2844), .ZN(n534) );
  LVT_AOI21HSV2 U2396 ( .A1(n2863), .A2(n534), .B(rw_P2_C2[1]), .ZN(n3075) );
  LVT_NAND2HSV2 U2397 ( .A1(n3075), .A2(rw_P2_C2[0]), .ZN(n2997) );
  LVT_NOR2HSV2 U2398 ( .A1(n2840), .A2(n2997), .ZN(n2775) );
  LVT_INOR2HSV1 U2399 ( .A1(debugStateC2[3]), .B1(debugStateC2[1]), .ZN(n2784)
         );
  LVT_CLKNHSV0 U2400 ( .I(debugStateC2[2]), .ZN(n2981) );
  LVT_INHSV2 U2401 ( .I(debugStateC2[0]), .ZN(n2785) );
  LVT_NAND3HSV2 U2402 ( .A1(n2784), .A2(n2981), .A3(n2785), .ZN(n693) );
  LVT_INHSV2 U2403 ( .I(n693), .ZN(n2955) );
  LVT_NAND2HSV2 U2404 ( .A1(n2775), .A2(n2955), .ZN(n2975) );
  LVT_INOR2HSV1 U2405 ( .A1(debugStateC2[1]), .B1(debugStateC2[0]), .ZN(n2980)
         );
  LVT_AND2HSV2 U2406 ( .A1(n2774), .A2(n2980), .Z(n1898) );
  LVT_CLKNHSV0 U2407 ( .I(n1898), .ZN(n2862) );
  LVT_AND2HSV2 U2408 ( .A1(n2975), .A2(n2862), .Z(n3039) );
  LVT_INHSV2 U2409 ( .I(n534), .ZN(n3099) );
  LVT_AOI21HSV2 U2410 ( .A1(n2775), .A2(n3070), .B(n3099), .ZN(n2776) );
  LVT_OA211HSV1 U2411 ( .A1(n2483), .A2(n420), .B(n3039), .C(n2776), .Z(n3032)
         );
  LVT_CLKNHSV0 U2412 ( .I(n3056), .ZN(n2860) );
  LVT_CLKNHSV0 U2413 ( .I(n3043), .ZN(n2960) );
  LVT_INHSV2 U2414 ( .I(n2959), .ZN(n2989) );
  LVT_NOR3HSV0 U2415 ( .A1(n2960), .A2(n2865), .A3(n2989), .ZN(n2777) );
  LVT_AOI211HSV0 U2416 ( .A1(n3060), .A2(n1674), .B(n3054), .C(n2777), .ZN(
        n2779) );
  LVT_OAI211HSV0 U2417 ( .A1(n2780), .A2(n2860), .B(n2779), .C(n2778), .ZN(
        n583) );
  LVT_CLKNHSV0 U2418 ( .I(n2011), .ZN(n2782) );
  LVT_NAND2HSV0 U2419 ( .A1(n3054), .A2(n3065), .ZN(n2781) );
  LVT_OAI211HSV1 U2420 ( .A1(n591), .A2(n592), .B(n2782), .C(n2781), .ZN(n464)
         );
  LVT_NOR2HSV0 U2421 ( .A1(n464), .A2(n465), .ZN(n463) );
  LVT_INOR2HSV1 U2422 ( .A1(n2784), .B1(n2783), .ZN(n3084) );
  LVT_CLKNAND2HSV0 U2423 ( .A1(n2784), .A2(debugStateC2[2]), .ZN(n2939) );
  LVT_INAND2HSV2 U2424 ( .A1(n2939), .B1(n2785), .ZN(n3006) );
  LVT_INAND2HSV2 U2425 ( .A1(n3084), .B1(n3006), .ZN(n500) );
  LVT_INAND2HSV2 U2426 ( .A1(n2939), .B1(debugStateC2[0]), .ZN(n2853) );
  LVT_INAND2HSV2 U2427 ( .A1(debugStateC2[3]), .B1(debugStateC2[2]), .ZN(n2938) );
  LVT_INAND2HSV2 U2428 ( .A1(n2938), .B1(n2980), .ZN(n2854) );
  LVT_NAND2HSV2 U2429 ( .A1(n2853), .A2(n2854), .ZN(n2861) );
  LVT_INHSV2 U2430 ( .I(n2938), .ZN(n2982) );
  LVT_NAND2HSV2 U2431 ( .A1(n2982), .A2(n2844), .ZN(n538) );
  LVT_INHSV2 U2432 ( .I(n538), .ZN(n3083) );
  LVT_XNOR2HSV1 U2433 ( .A1(addr_C2_M[9]), .A2(addr_P2_C2[9]), .ZN(n2789) );
  LVT_XNOR2HSV1 U2434 ( .A1(addr_C2_M[11]), .A2(addr_P2_C2[11]), .ZN(n2788) );
  LVT_XNOR2HSV1 U2435 ( .A1(addr_C2_M[5]), .A2(addr_P2_C2[5]), .ZN(n2787) );
  LVT_XNOR2HSV0 U2436 ( .A1(addr_C2_M[12]), .A2(addr_P2_C2[12]), .ZN(n2786) );
  LVT_NAND4HSV2 U2437 ( .A1(n2789), .A2(n2788), .A3(n2787), .A4(n2786), .ZN(
        n2795) );
  LVT_XNOR2HSV1 U2438 ( .A1(addr_C2_M[1]), .A2(addr_P2_C2[1]), .ZN(n2793) );
  LVT_XNOR2HSV1 U2439 ( .A1(addr_C2_M[6]), .A2(addr_P2_C2[6]), .ZN(n2792) );
  LVT_XNOR2HSV1 U2440 ( .A1(addr_C2_M[3]), .A2(n1290), .ZN(n2791) );
  LVT_XNOR2HSV1 U2441 ( .A1(addr_C2_M[15]), .A2(addr_P2_C2[15]), .ZN(n2790) );
  LVT_NAND4HSV2 U2442 ( .A1(n2793), .A2(n2792), .A3(n2791), .A4(n2790), .ZN(
        n2794) );
  LVT_NOR2HSV2 U2443 ( .A1(n2795), .A2(n2794), .ZN(n2807) );
  LVT_XNOR2HSV1 U2444 ( .A1(addr_C2_M[14]), .A2(addr_P2_C2[14]), .ZN(n2799) );
  LVT_XNOR2HSV1 U2445 ( .A1(addr_C2_M[10]), .A2(addr_P2_C2[10]), .ZN(n2798) );
  LVT_XNOR2HSV1 U2446 ( .A1(addr_C2_M[13]), .A2(addr_P2_C2[13]), .ZN(n2797) );
  LVT_XNOR2HSV1 U2447 ( .A1(addr_C2_M[8]), .A2(addr_P2_C2[8]), .ZN(n2796) );
  LVT_NAND4HSV2 U2448 ( .A1(n2799), .A2(n2798), .A3(n2797), .A4(n2796), .ZN(
        n2805) );
  LVT_INHSV2 U2449 ( .I(addr_P2_C2[0]), .ZN(n3092) );
  LVT_XOR2HSV0 U2450 ( .A1(addr_C2_M[0]), .A2(n3092), .Z(n2803) );
  LVT_XNOR2HSV1 U2451 ( .A1(addr_C2_M[7]), .A2(addr_P2_C2[7]), .ZN(n2802) );
  LVT_XNOR2HSV1 U2452 ( .A1(addr_C2_M[2]), .A2(addr_P2_C2[2]), .ZN(n2801) );
  LVT_XNOR2HSV1 U2453 ( .A1(addr_C2_M[4]), .A2(addr_P2_C2[4]), .ZN(n2800) );
  LVT_NAND4HSV2 U2454 ( .A1(n2803), .A2(n2802), .A3(n2801), .A4(n2800), .ZN(
        n2804) );
  LVT_NOR2HSV2 U2455 ( .A1(n2805), .A2(n2804), .ZN(n2806) );
  LVT_NAND2HSV2 U2456 ( .A1(n2807), .A2(n2806), .ZN(n2808) );
  LVT_NAND2HSV2 U2457 ( .A1(n2809), .A2(n2808), .ZN(n2852) );
  LVT_NAND2HSV2 U2458 ( .A1(n2852), .A2(en_M_C2), .ZN(n3004) );
  LVT_INHSV2 U2459 ( .I(n2809), .ZN(n2846) );
  LVT_OR2HSV1 U2460 ( .A1(n3004), .A2(n2846), .Z(n2952) );
  LVT_INHSV2 U2461 ( .I(n2952), .ZN(n3029) );
  LVT_NOR2HSV1 U2462 ( .A1(n3004), .A2(n538), .ZN(n3071) );
  LVT_XNOR2HSV0 U2463 ( .A1(allowReadAddr_C1_C2[1]), .A2(addr_P1_C1[1]), .ZN(
        n2812) );
  LVT_XNOR2HSV0 U2464 ( .A1(allowReadAddr_C1_C2[7]), .A2(addr_P1_C1[7]), .ZN(
        n2811) );
  LVT_NAND3HSV2 U2465 ( .A1(n2812), .A2(n2811), .A3(n2810), .ZN(n2815) );
  LVT_XOR2HSV0 U2466 ( .A1(allowReadAddr_C1_C2[0]), .A2(addr_P1_C1[0]), .Z(
        n2814) );
  LVT_XOR2HSV0 U2467 ( .A1(allowReadAddr_C1_C2[2]), .A2(addr_P1_C1[2]), .Z(
        n2813) );
  LVT_NOR3HSV2 U2468 ( .A1(n2815), .A2(n2814), .A3(n2813), .ZN(n2832) );
  LVT_XNOR2HSV0 U2469 ( .A1(allowReadAddr_C1_C2[8]), .A2(addr_P1_C1[8]), .ZN(
        n2819) );
  LVT_XNOR2HSV0 U2470 ( .A1(allowReadAddr_C1_C2[14]), .A2(addr_P1_C1[14]), 
        .ZN(n2818) );
  LVT_XNOR2HSV0 U2471 ( .A1(allowReadAddr_C1_C2[11]), .A2(addr_P1_C1[11]), 
        .ZN(n2817) );
  LVT_XNOR2HSV0 U2472 ( .A1(allowReadAddr_C1_C2[4]), .A2(addr_P1_C1[4]), .ZN(
        n2816) );
  LVT_NAND4HSV2 U2473 ( .A1(n2819), .A2(n2818), .A3(n2817), .A4(n2816), .ZN(
        n2825) );
  LVT_XNOR2HSV0 U2474 ( .A1(allowReadAddr_C1_C2[6]), .A2(addr_P1_C1[6]), .ZN(
        n2823) );
  LVT_XNOR2HSV0 U2475 ( .A1(allowReadAddr_C1_C2[10]), .A2(addr_P1_C1[10]), 
        .ZN(n2822) );
  LVT_XNOR2HSV0 U2476 ( .A1(allowReadAddr_C1_C2[13]), .A2(addr_P1_C1[13]), 
        .ZN(n2821) );
  LVT_XNOR2HSV0 U2477 ( .A1(allowReadAddr_C1_C2[15]), .A2(addr_P1_C1[15]), 
        .ZN(n2820) );
  LVT_NAND4HSV2 U2478 ( .A1(n2823), .A2(n2822), .A3(n2821), .A4(n2820), .ZN(
        n2824) );
  LVT_NOR2HSV2 U2479 ( .A1(n2825), .A2(n2824), .ZN(n2831) );
  LVT_XNOR2HSV0 U2480 ( .A1(allowReadAddr_C1_C2[5]), .A2(addr_P1_C1[5]), .ZN(
        n2829) );
  LVT_XNOR2HSV0 U2481 ( .A1(allowReadAddr_C1_C2[9]), .A2(addr_P1_C1[9]), .ZN(
        n2828) );
  LVT_XNOR2HSV0 U2482 ( .A1(allowReadAddr_C1_C2[12]), .A2(addr_P1_C1[12]), 
        .ZN(n2827) );
  LVT_XNOR2HSV0 U2483 ( .A1(allowReadAddr_C1_C2[3]), .A2(addr_P1_C1[3]), .ZN(
        n2826) );
  LVT_AND4HSV1 U2484 ( .A1(n2829), .A2(n2828), .A3(n2827), .A4(n2826), .Z(
        n2830) );
  LVT_NAND3HSV2 U2485 ( .A1(n2832), .A2(n2831), .A3(n2830), .ZN(n1555) );
  LVT_INHSV2 U2486 ( .I(n1555), .ZN(n2924) );
  LVT_NOR2HSV2 U2487 ( .A1(n2833), .A2(n2924), .ZN(n2968) );
  LVT_INAND2HSV2 U2488 ( .A1(n2959), .B1(n3068), .ZN(n2964) );
  LVT_CLKNHSV0 U2489 ( .I(en_M_C1), .ZN(n3064) );
  LVT_NOR2HSV0 U2490 ( .A1(n1674), .A2(n639), .ZN(n3036) );
  LVT_NOR2HSV0 U2491 ( .A1(rw_P1_C1[1]), .A2(rw_P1_C1[0]), .ZN(n2857) );
  LVT_IOA21HSV2 U2492 ( .A1(n2958), .A2(n2857), .B(n2959), .ZN(n2838) );
  LVT_CLKNHSV0 U2493 ( .I(n2835), .ZN(n2836) );
  LVT_AOI21HSV0 U2494 ( .A1(n2987), .A2(n2836), .B(en_M_C1), .ZN(n2837) );
  LVT_AOI211HSV0 U2495 ( .A1(n3055), .A2(n2838), .B(n2837), .C(n3036), .ZN(
        n932) );
  LVT_AND2HSV2 U2496 ( .A1(n3075), .A2(n3076), .Z(n3074) );
  LVT_INAND3HSV2 U2497 ( .A1(n2840), .B1(n3070), .B2(n3074), .ZN(n3025) );
  LVT_CLKNHSV0 U2498 ( .I(n3025), .ZN(n2839) );
  LVT_AOI211HSV0 U2499 ( .A1(n3084), .A2(n3004), .B(n3099), .C(n2839), .ZN(
        n2842) );
  LVT_INAND2HSV2 U2500 ( .A1(n2840), .B1(n2955), .ZN(n2956) );
  LVT_INHSV2 U2501 ( .I(n3074), .ZN(n3000) );
  LVT_NOR2HSV2 U2502 ( .A1(n2956), .A2(n3000), .ZN(n3073) );
  LVT_INHSV2 U2503 ( .I(n3073), .ZN(n2841) );
  LVT_OAI211HSV0 U2504 ( .A1(n2843), .A2(n420), .B(n2842), .C(n2841), .ZN(n685) );
  LVT_NOR2HSV0 U2505 ( .A1(debugStateC2[2]), .A2(debugStateC2[3]), .ZN(n2845)
         );
  LVT_NAND2HSV2 U2506 ( .A1(n2845), .A2(n2844), .ZN(n1849) );
  LVT_CLKNHSV0 U2507 ( .I(rw_C2_M[1]), .ZN(n2944) );
  LVT_OAI211HSV0 U2508 ( .A1(n420), .A2(n2944), .B(n2846), .C(n1849), .ZN(n418) );
  LVT_AND2HSV2 U2509 ( .A1(n2845), .A2(n2980), .Z(n3046) );
  LVT_NAND2HSV0 U2510 ( .A1(n3046), .A2(en_M_C2), .ZN(n1780) );
  LVT_NAND2HSV0 U2511 ( .A1(n1780), .A2(n1849), .ZN(n1901) );
  LVT_CLKNHSV0 U2512 ( .I(n1901), .ZN(n2848) );
  LVT_NAND3HSV2 U2513 ( .A1(n3078), .A2(n3070), .A3(n3077), .ZN(n417) );
  LVT_OAI211HSV0 U2514 ( .A1(n2848), .A2(n2847), .B(n417), .C(n2846), .ZN(
        n2851) );
  LVT_INAND3HSV2 U2515 ( .A1(n2849), .B1(n2955), .B2(n3077), .ZN(n513) );
  LVT_CLKNHSV0 U2516 ( .I(n513), .ZN(n2850) );
  LVT_AOI211HSV0 U2517 ( .A1(n3047), .A2(en_C2_P2), .B(n2851), .C(n2850), .ZN(
        n574) );
  LVT_NAND2HSV0 U2518 ( .A1(n2926), .A2(n2855), .ZN(n2928) );
  LVT_NOR2HSV1 U2519 ( .A1(n1672), .A2(C1_stall), .ZN(n2856) );
  LVT_CLKNAND2HSV1 U2520 ( .A1(n2929), .A2(n2856), .ZN(n2966) );
  LVT_AND2HSV2 U2521 ( .A1(n3054), .A2(n2857), .Z(n3044) );
  LVT_CLKNHSV1 U2522 ( .I(rw_C1_M[1]), .ZN(n2937) );
  LVT_INHSV2 U2523 ( .I(n1789), .ZN(n2950) );
  LVT_OAI211HSV0 U2524 ( .A1(n2860), .A2(n2937), .B(n2950), .C(n600), .ZN(n716) );
  LVT_INOR2HSV0 U2525 ( .A1(n2861), .B1(n3004), .ZN(n2394) );
  LVT_AOI21HSV0 U2526 ( .A1(n3006), .A2(n2862), .B(n3004), .ZN(n691) );
  LVT_NAND2HSV2 U2527 ( .A1(n694), .A2(n3003), .ZN(n440) );
  HVT_AOI21HSV0 U2528 ( .A1(n3003), .A2(n3078), .B(n444), .ZN(n3035) );
  LVT_CLKNHSV0 U2529 ( .I(n3035), .ZN(n1274) );
  LVT_INOR2HSV1 U2530 ( .A1(n2864), .B1(n2969), .ZN(n641) );
  LVT_CLKNHSV0 U2531 ( .I(n3053), .ZN(n2866) );
  LVT_AOI21HSV2 U2532 ( .A1(n2866), .A2(n2959), .B(n2865), .ZN(n2407) );
  LVT_CLKNHSV1 U2533 ( .I(n2407), .ZN(n1624) );
  LVT_CLKNHSV0 U2534 ( .I(pc_proc1_code1[7]), .ZN(n2867) );
  LVT_CLKNHSV0 U2535 ( .I(pc_proc1_code1[0]), .ZN(P1_N104) );
  LVT_CLKNHSV0 U2536 ( .I(pc_proc1_code1[1]), .ZN(n2946) );
  LVT_INOR3HSV2 U2537 ( .A1(pc_proc1_code1[2]), .B1(P1_N104), .B2(n2946), .ZN(
        n2991) );
  LVT_NAND2HSV0 U2538 ( .A1(n2991), .A2(pc_proc1_code1[3]), .ZN(n2990) );
  LVT_CLKNHSV0 U2539 ( .I(pc_proc1_code1[4]), .ZN(n2936) );
  LVT_NOR2HSV2 U2540 ( .A1(n2990), .A2(n2936), .ZN(n2935) );
  LVT_INHSV2 U2541 ( .I(n2935), .ZN(n2917) );
  LVT_CLKNHSV0 U2542 ( .I(pc_proc1_code1[5]), .ZN(n2916) );
  LVT_NOR2HSV2 U2543 ( .A1(n2917), .A2(n2916), .ZN(n3012) );
  LVT_NAND2HSV0 U2544 ( .A1(n3012), .A2(pc_proc1_code1[6]), .ZN(n3011) );
  LVT_MUX2NHSV0 U2545 ( .I0(pc_proc1_code1[7]), .I1(n2867), .S(n3011), .ZN(
        P1_N111) );
  LVT_CLKNHSV0 U2546 ( .I(pc_proc2_code2[7]), .ZN(n2868) );
  LVT_CLKNHSV0 U2547 ( .I(pc_proc2_code2[0]), .ZN(P2_N104) );
  LVT_CLKNHSV0 U2548 ( .I(pc_proc2_code2[1]), .ZN(n2942) );
  LVT_INOR3HSV2 U2549 ( .A1(pc_proc2_code2[2]), .B1(P2_N104), .B2(n2942), .ZN(
        n2993) );
  LVT_NAND2HSV0 U2550 ( .A1(n2993), .A2(pc_proc2_code2[3]), .ZN(n2992) );
  LVT_CLKNHSV0 U2551 ( .I(pc_proc2_code2[4]), .ZN(n2934) );
  LVT_NOR2HSV2 U2552 ( .A1(n2992), .A2(n2934), .ZN(n2933) );
  LVT_INHSV2 U2553 ( .I(n2933), .ZN(n2922) );
  LVT_CLKNHSV0 U2554 ( .I(pc_proc2_code2[5]), .ZN(n2921) );
  LVT_NOR2HSV2 U2555 ( .A1(n2922), .A2(n2921), .ZN(n3014) );
  LVT_NAND2HSV0 U2556 ( .A1(n3014), .A2(pc_proc2_code2[6]), .ZN(n3013) );
  LVT_MUX2NHSV0 U2557 ( .I0(pc_proc2_code2[7]), .I1(n2868), .S(n3013), .ZN(
        P2_N111) );
  LVT_XOR2HSV0 U2558 ( .A1(allowReadAddr_C1_C2[0]), .A2(n3092), .Z(n2870) );
  LVT_INHSV2 U2559 ( .I(allowRead_C1_C2), .ZN(n2906) );
  LVT_XNOR2HSV1 U2560 ( .A1(allowReadAddr_C1_C2[14]), .A2(addr_P2_C2[14]), 
        .ZN(n2869) );
  LVT_NAND3HSV2 U2561 ( .A1(n2870), .A2(n2906), .A3(n2869), .ZN(n2873) );
  LVT_XOR2HSV0 U2562 ( .A1(allowReadAddr_C1_C2[2]), .A2(addr_P2_C2[2]), .Z(
        n2872) );
  LVT_XOR2HSV0 U2563 ( .A1(allowReadAddr_C1_C2[3]), .A2(n1290), .Z(n2871) );
  LVT_NOR3HSV2 U2564 ( .A1(n2873), .A2(n2872), .A3(n2871), .ZN(n2890) );
  LVT_XNOR2HSV1 U2565 ( .A1(allowReadAddr_C1_C2[9]), .A2(addr_P2_C2[9]), .ZN(
        n2877) );
  LVT_XNOR2HSV1 U2566 ( .A1(allowReadAddr_C1_C2[1]), .A2(addr_P2_C2[1]), .ZN(
        n2876) );
  LVT_XNOR2HSV1 U2567 ( .A1(allowReadAddr_C1_C2[5]), .A2(addr_P2_C2[5]), .ZN(
        n2875) );
  LVT_XNOR2HSV1 U2568 ( .A1(allowReadAddr_C1_C2[10]), .A2(addr_P2_C2[10]), 
        .ZN(n2874) );
  LVT_AND4HSV1 U2569 ( .A1(n2877), .A2(n2876), .A3(n2875), .A4(n2874), .Z(
        n2889) );
  LVT_XNOR2HSV1 U2570 ( .A1(allowReadAddr_C1_C2[7]), .A2(addr_P2_C2[7]), .ZN(
        n2881) );
  LVT_XNOR2HSV1 U2571 ( .A1(allowReadAddr_C1_C2[11]), .A2(addr_P2_C2[11]), 
        .ZN(n2880) );
  LVT_XNOR2HSV1 U2572 ( .A1(allowReadAddr_C1_C2[8]), .A2(addr_P2_C2[8]), .ZN(
        n2879) );
  LVT_XNOR2HSV1 U2573 ( .A1(allowReadAddr_C1_C2[13]), .A2(addr_P2_C2[13]), 
        .ZN(n2878) );
  LVT_NAND4HSV2 U2574 ( .A1(n2881), .A2(n2880), .A3(n2879), .A4(n2878), .ZN(
        n2887) );
  LVT_XNOR2HSV1 U2575 ( .A1(allowReadAddr_C1_C2[6]), .A2(addr_P2_C2[6]), .ZN(
        n2885) );
  LVT_XNOR2HSV1 U2576 ( .A1(allowReadAddr_C1_C2[15]), .A2(addr_P2_C2[15]), 
        .ZN(n2884) );
  LVT_XNOR2HSV1 U2577 ( .A1(allowReadAddr_C1_C2[4]), .A2(addr_P2_C2[4]), .ZN(
        n2883) );
  LVT_XNOR2HSV0 U2578 ( .A1(allowReadAddr_C1_C2[12]), .A2(addr_P2_C2[12]), 
        .ZN(n2882) );
  LVT_NAND4HSV2 U2579 ( .A1(n2885), .A2(n2884), .A3(n2883), .A4(n2882), .ZN(
        n2886) );
  LVT_NOR2HSV2 U2580 ( .A1(n2887), .A2(n2886), .ZN(n2888) );
  LVT_NAND3HSV2 U2581 ( .A1(n2890), .A2(n2889), .A3(n2888), .ZN(n3015) );
  LVT_CLKNHSV0 U2582 ( .I(n2997), .ZN(n2915) );
  LVT_XNOR2HSV1 U2583 ( .A1(allowReadAddr_C2_C1[6]), .A2(addr_P2_C2[6]), .ZN(
        n2894) );
  LVT_XNOR2HSV1 U2584 ( .A1(allowReadAddr_C2_C1[5]), .A2(addr_P2_C2[5]), .ZN(
        n2893) );
  LVT_XNOR2HSV1 U2585 ( .A1(allowReadAddr_C2_C1[9]), .A2(addr_P2_C2[9]), .ZN(
        n2892) );
  LVT_XNOR2HSV1 U2586 ( .A1(allowReadAddr_C2_C1[1]), .A2(addr_P2_C2[1]), .ZN(
        n2891) );
  LVT_NAND4HSV2 U2587 ( .A1(n2894), .A2(n2893), .A3(n2892), .A4(n2891), .ZN(
        n2900) );
  LVT_XNOR2HSV1 U2588 ( .A1(allowReadAddr_C2_C1[3]), .A2(n1290), .ZN(n2898) );
  LVT_XNOR2HSV1 U2589 ( .A1(allowReadAddr_C2_C1[14]), .A2(addr_P2_C2[14]), 
        .ZN(n2897) );
  LVT_XNOR2HSV1 U2590 ( .A1(allowReadAddr_C2_C1[4]), .A2(addr_P2_C2[4]), .ZN(
        n2896) );
  LVT_XNOR2HSV1 U2591 ( .A1(allowReadAddr_C2_C1[10]), .A2(addr_P2_C2[10]), 
        .ZN(n2895) );
  LVT_NAND4HSV2 U2592 ( .A1(n2898), .A2(n2897), .A3(n2896), .A4(n2895), .ZN(
        n2899) );
  LVT_NOR2HSV2 U2593 ( .A1(n2900), .A2(n2899), .ZN(n2914) );
  LVT_XNOR2HSV1 U2594 ( .A1(allowReadAddr_C2_C1[2]), .A2(addr_P2_C2[2]), .ZN(
        n2904) );
  LVT_XNOR2HSV1 U2595 ( .A1(allowReadAddr_C2_C1[11]), .A2(addr_P2_C2[11]), 
        .ZN(n2903) );
  LVT_XNOR2HSV1 U2596 ( .A1(allowReadAddr_C2_C1[13]), .A2(addr_P2_C2[13]), 
        .ZN(n2902) );
  LVT_XNOR2HSV0 U2597 ( .A1(allowReadAddr_C2_C1[0]), .A2(addr_P2_C2[0]), .ZN(
        n2901) );
  LVT_AND4HSV1 U2598 ( .A1(n2904), .A2(n2903), .A3(n2902), .A4(n2901), .Z(
        n2913) );
  LVT_XNOR2HSV1 U2599 ( .A1(allowReadAddr_C2_C1[15]), .A2(addr_P2_C2[15]), 
        .ZN(n2907) );
  LVT_XNOR2HSV1 U2600 ( .A1(allowReadAddr_C2_C1[7]), .A2(addr_P2_C2[7]), .ZN(
        n2905) );
  LVT_NAND3HSV2 U2601 ( .A1(n2907), .A2(n2906), .A3(n2905), .ZN(n2911) );
  LVT_XNOR2HSV1 U2602 ( .A1(allowReadAddr_C2_C1[8]), .A2(addr_P2_C2[8]), .ZN(
        n2909) );
  LVT_XNOR2HSV0 U2603 ( .A1(allowReadAddr_C2_C1[12]), .A2(addr_P2_C2[12]), 
        .ZN(n2908) );
  LVT_NAND2HSV2 U2604 ( .A1(n2909), .A2(n2908), .ZN(n2910) );
  LVT_NOR2HSV2 U2605 ( .A1(n2911), .A2(n2910), .ZN(n2912) );
  LVT_NAND3HSV2 U2606 ( .A1(n2914), .A2(n2913), .A3(n2912), .ZN(n2923) );
  LVT_OAI22HSV0 U2607 ( .A1(n3074), .A2(n3015), .B1(n2915), .B2(n2923), .ZN(
        n1740) );
  LVT_AOI21HSV1 U2608 ( .A1(n2917), .A2(n2916), .B(n3012), .ZN(P1_N109) );
  LVT_NAND3HSV0 U2609 ( .A1(n2923), .A2(en_M_C2), .A3(n3037), .ZN(n2920) );
  HVT_NOR2HSV0 U2610 ( .A1(debugStateC2[1]), .A2(debugStateC2[0]), .ZN(n2918)
         );
  LVT_CLKNAND2HSV1 U2611 ( .A1(n2982), .A2(n2918), .ZN(n3027) );
  LVT_INHSV2 U2612 ( .I(en_M_C2), .ZN(n3098) );
  LVT_NOR2HSV2 U2613 ( .A1(n3027), .A2(n3098), .ZN(n2919) );
  LVT_NAND2HSV2 U2614 ( .A1(n3015), .A2(n2919), .ZN(n2953) );
  LVT_CLKNAND2HSV1 U2615 ( .A1(n2920), .A2(n2953), .ZN(n536) );
  LVT_AOI21HSV1 U2616 ( .A1(n2922), .A2(n2921), .B(n3014), .ZN(P2_N109) );
  LVT_INHSV2 U2617 ( .I(n2923), .ZN(n2999) );
  LVT_AOI21HSV0 U2618 ( .A1(n3074), .A2(n2999), .B(n3072), .ZN(n537) );
  LVT_NAND2HSV0 U2619 ( .A1(n2924), .A2(n3066), .ZN(n2925) );
  LVT_OAI211HSV0 U2620 ( .A1(n3066), .A2(n2929), .B(n3053), .C(n2925), .ZN(
        n1543) );
  LVT_CLKNHSV0 U2621 ( .I(n3075), .ZN(n2391) );
  LVT_NAND3HSV2 U2622 ( .A1(n1555), .A2(en_M_C1), .A3(n3041), .ZN(n2972) );
  LVT_NOR2HSV1 U2623 ( .A1(n2928), .A2(debugStateC1[0]), .ZN(n3049) );
  LVT_NAND2HSV0 U2624 ( .A1(n2972), .A2(n2965), .ZN(n1791) );
  LVT_NOR2HSV1 U2625 ( .A1(n2931), .A2(n2930), .ZN(n3045) );
  LVT_CLKNHSV0 U2626 ( .I(n3069), .ZN(n1819) );
  LVT_NAND2HSV0 U2627 ( .A1(n2987), .A2(n2932), .ZN(n1804) );
  LVT_AOI21HSV0 U2628 ( .A1(n2992), .A2(n2934), .B(n2933), .ZN(P2_N108) );
  LVT_AOI21HSV0 U2629 ( .A1(n2990), .A2(n2936), .B(n2935), .ZN(P1_N108) );
  LVT_CLKNHSV0 U2630 ( .I(n600), .ZN(n2570) );
  LVT_INHSV2 U2631 ( .I(mb_prefer), .ZN(n2452) );
  LVT_OR2HSV1 U2632 ( .A1(rw_C1_M[0]), .A2(n2937), .Z(n711) );
  LVT_NAND2HSV2 U2633 ( .A1(n2452), .A2(n711), .ZN(n707) );
  LVT_CLKNHSV0 U2634 ( .I(rw_C2_M[0]), .ZN(n2943) );
  LVT_NAND2HSV2 U2635 ( .A1(rw_C2_M[1]), .A2(n2943), .ZN(n712) );
  LVT_AOI21HSV0 U2636 ( .A1(n707), .A2(n712), .B(n2937), .ZN(n709) );
  LVT_CLKNHSV0 U2637 ( .I(n3044), .ZN(n1801) );
  HVT_CLKNHSV0 U2638 ( .I(debugStateC2[1]), .ZN(n2941) );
  LVT_OAI21HSV0 U2639 ( .A1(n2939), .A2(en_M_C2), .B(n2938), .ZN(n2940) );
  LVT_OAI21HSV0 U2640 ( .A1(n3098), .A2(n2941), .B(n2940), .ZN(n543) );
  LVT_AND2HSV2 U2641 ( .A1(n3054), .A2(C1_stall), .Z(n3038) );
  LVT_CLKNHSV0 U2642 ( .I(n3038), .ZN(n1553) );
  LVT_CLKNHSV0 U2643 ( .I(n639), .ZN(n3062) );
  LVT_NOR2HSV1 U2644 ( .A1(P2_N104), .A2(n2942), .ZN(n2977) );
  LVT_AOI21HSV0 U2645 ( .A1(P2_N104), .A2(n2942), .B(n2977), .ZN(P2_N105) );
  LVT_OAI32HSV0 U2646 ( .A1(n2944), .A2(n2943), .A3(n2452), .B1(n711), .B2(
        n2944), .ZN(n710) );
  LVT_NOR3HSV2 U2647 ( .A1(debugDelay[2]), .A2(debugDelay[1]), .A3(
        debugDelay[0]), .ZN(n2451) );
  LVT_CLKNHSV0 U2648 ( .I(n2451), .ZN(n1442) );
  LVT_NOR2HSV1 U2649 ( .A1(debugDelay[1]), .A2(debugDelay[0]), .ZN(n2947) );
  LVT_CLKNHSV0 U2650 ( .I(debugDelay[2]), .ZN(n2945) );
  LVT_OAI21HSV0 U2651 ( .A1(n2947), .A2(n2945), .B(n1442), .ZN(n1441) );
  LVT_NOR2HSV1 U2652 ( .A1(P1_N104), .A2(n2946), .ZN(n2978) );
  LVT_AOI21HSV0 U2653 ( .A1(P1_N104), .A2(n2946), .B(n2978), .ZN(P1_N105) );
  LVT_INHSV2 U2654 ( .I(ins_code2_proc2[20]), .ZN(n2587) );
  LVT_INHSV2 U2655 ( .I(ins_code2_proc2[21]), .ZN(n2586) );
  LVT_OAI22HSV2 U2656 ( .A1(n2587), .A2(n2586), .B1(ins_code2_proc2[21]), .B2(
        ins_code2_proc2[20]), .ZN(n2948) );
  LVT_NOR2HSV2 U2657 ( .A1(n2948), .A2(ins_code2_proc2[22]), .ZN(n548) );
  LVT_CLKNHSV0 U2658 ( .I(ins_code2_proc2[23]), .ZN(n2582) );
  LVT_NAND3HSV1 U2659 ( .A1(en_C2_P2), .A2(n548), .A3(n2582), .ZN(n554) );
  LVT_INHSV2 U2660 ( .I(ins_code1_proc1[20]), .ZN(n2592) );
  LVT_INHSV2 U2661 ( .I(ins_code1_proc1[21]), .ZN(n2591) );
  LVT_OAI22HSV2 U2662 ( .A1(n2592), .A2(n2591), .B1(ins_code1_proc1[21]), .B2(
        ins_code1_proc1[20]), .ZN(n2949) );
  LVT_NOR2HSV2 U2663 ( .A1(n2949), .A2(ins_code1_proc1[22]), .ZN(n650) );
  LVT_CLKNHSV0 U2664 ( .I(ins_code1_proc1[23]), .ZN(n2588) );
  LVT_NAND3HSV1 U2665 ( .A1(n650), .A2(en_C1_P1), .A3(n2588), .ZN(n656) );
  LVT_AO21HSV0 U2666 ( .A1(debugDelay[0]), .A2(debugDelay[1]), .B(n2947), .Z(
        n1438) );
  LVT_NOR2HSV0 U2667 ( .A1(ins_code1_proc1[20]), .A2(ins_code1_proc1[21]), 
        .ZN(n662) );
  LVT_CLKNHSV0 U2668 ( .I(ins_code1_proc1[22]), .ZN(n2590) );
  LVT_OAI21HSV1 U2669 ( .A1(n662), .A2(n2590), .B(n2949), .ZN(n655) );
  LVT_NOR2HSV0 U2670 ( .A1(ins_code2_proc2[20]), .A2(ins_code2_proc2[21]), 
        .ZN(n560) );
  LVT_CLKNHSV0 U2671 ( .I(ins_code2_proc2[22]), .ZN(n2584) );
  LVT_OAI21HSV1 U2672 ( .A1(n560), .A2(n2584), .B(n2948), .ZN(n553) );
  LVT_NOR3HSV1 U2673 ( .A1(n2586), .A2(ins_code2_proc2[22]), .A3(
        ins_code2_proc2[20]), .ZN(n564) );
  LVT_CLKNHSV0 U2674 ( .I(n564), .ZN(n2585) );
  LVT_CLKNHSV0 U2675 ( .I(n2948), .ZN(n565) );
  LVT_AOI21HSV0 U2676 ( .A1(ins_code2_proc2[20]), .A2(n2586), .B(n564), .ZN(
        n570) );
  LVT_CLKNHSV0 U2677 ( .I(n2949), .ZN(n667) );
  LVT_NOR3HSV1 U2678 ( .A1(ins_code1_proc1[22]), .A2(ins_code1_proc1[20]), 
        .A3(n2591), .ZN(n666) );
  LVT_AOI21HSV0 U2679 ( .A1(ins_code1_proc1[20]), .A2(n2591), .B(n666), .ZN(
        n672) );
  LVT_CLKNHSV1 U2680 ( .I(allowReadAddr_C2_C1[6]), .ZN(n2479) );
  LVT_CLKNHSV0 U2681 ( .I(addr_C2_M[0]), .ZN(n2437) );
  LVT_CLKNHSV1 U2682 ( .I(allowReadAddr_C2_C1[4]), .ZN(n2478) );
  LVT_CLKNHSV0 U2683 ( .I(addr_C2_M[6]), .ZN(n2443) );
  LVT_CLKNHSV0 U2684 ( .I(addr_C2_C1[0]), .ZN(n2438) );
  LVT_CLKNHSV0 U2685 ( .I(addr_C2_M[12]), .ZN(n2450) );
  LVT_CLKNHSV0 U2686 ( .I(addr_C2_M[10]), .ZN(n2441) );
  LVT_CLKNHSV0 U2687 ( .I(addr_C2_M[9]), .ZN(n2447) );
  LVT_CLKNHSV0 U2688 ( .I(addr_C2_M[5]), .ZN(n2448) );
  LVT_CLKNHSV1 U2689 ( .I(allowReadAddr_C1_C2[15]), .ZN(n2486) );
  LVT_CLKNHSV0 U2690 ( .I(addr_C2_M[2]), .ZN(n2427) );
  LVT_CLKNHSV0 U2691 ( .I(addr_C2_M[1]), .ZN(n2416) );
  LVT_CLKNHSV1 U2692 ( .I(addr_P1_C1[15]), .ZN(n2577) );
  LVT_CLKNHSV0 U2693 ( .I(allowReadAddr_C1_C2[1]), .ZN(n2507) );
  LVT_CLKNHSV1 U2694 ( .I(addr_P1_C1[1]), .ZN(n2551) );
  LVT_CLKNHSV0 U2695 ( .I(allowReadAddr_C1_C2[2]), .ZN(n2506) );
  LVT_CLKNHSV0 U2696 ( .I(allowReadAddr_C2_C1[13]), .ZN(n2505) );
  LVT_CLKNHSV0 U2697 ( .I(allowReadAddr_C2_C1[14]), .ZN(n2504) );
  LVT_CLKNHSV0 U2698 ( .I(allowReadAddr_C2_C1[15]), .ZN(n2503) );
  LVT_CLKNHSV0 U2699 ( .I(addr_P1_C1[2]), .ZN(n2549) );
  LVT_CLKNHSV0 U2700 ( .I(addr_C2_M[15]), .ZN(n2439) );
  LVT_CLKNHSV0 U2701 ( .I(allowReadAddr_C1_C2[3]), .ZN(n2502) );
  LVT_CLKNHSV1 U2702 ( .I(addr_P1_C1[14]), .ZN(n2509) );
  LVT_CLKNHSV1 U2703 ( .I(addr_P1_C1[3]), .ZN(n2581) );
  LVT_CLKNHSV1 U2704 ( .I(allowReadAddr_C1_C2[4]), .ZN(n2480) );
  LVT_CLKNHSV0 U2705 ( .I(addr_C2_M[8]), .ZN(n2440) );
  LVT_CLKNHSV0 U2706 ( .I(addr_C1_M[5]), .ZN(n2433) );
  LVT_CLKNHSV0 U2707 ( .I(addr_C1_M[6]), .ZN(n2432) );
  LVT_CLKNHSV0 U2708 ( .I(addr_C1_M[7]), .ZN(n2431) );
  LVT_CLKNHSV0 U2709 ( .I(addr_C1_M[9]), .ZN(n2430) );
  LVT_CLKNHSV0 U2710 ( .I(addr_C1_M[10]), .ZN(n2429) );
  LVT_CLKNHSV0 U2711 ( .I(addr_C1_M[11]), .ZN(n2428) );
  LVT_CLKNHSV0 U2712 ( .I(addr_C2_M[3]), .ZN(n2426) );
  LVT_CLKNHSV0 U2713 ( .I(addr_C1_M[15]), .ZN(n2425) );
  LVT_CLKNHSV0 U2714 ( .I(addr_C2_C1[4]), .ZN(n2457) );
  LVT_CLKNHSV0 U2715 ( .I(addr_C2_C1[8]), .ZN(n2458) );
  LVT_CLKNHSV0 U2716 ( .I(addr_C1_M[1]), .ZN(n2424) );
  LVT_CLKNHSV0 U2717 ( .I(addr_C2_C1[15]), .ZN(n2459) );
  LVT_CLKNHSV0 U2718 ( .I(addr_C1_M[2]), .ZN(n2423) );
  LVT_CLKNHSV1 U2719 ( .I(addr_C2_C1[3]), .ZN(n2460) );
  LVT_CLKNHSV0 U2720 ( .I(addr_C1_M[3]), .ZN(n2422) );
  LVT_CLKNHSV0 U2721 ( .I(addr_C2_C1[2]), .ZN(n2461) );
  LVT_CLKNHSV0 U2722 ( .I(addr_C1_M[4]), .ZN(n2421) );
  LVT_CLKNHSV0 U2723 ( .I(addr_C2_C1[1]), .ZN(n2462) );
  LVT_CLKNHSV0 U2724 ( .I(addr_C1_M[8]), .ZN(n2420) );
  LVT_CLKNHSV0 U2725 ( .I(addr_C1_M[12]), .ZN(n2419) );
  LVT_CLKNHSV0 U2726 ( .I(addr_C1_M[13]), .ZN(n2418) );
  LVT_CLKNHSV0 U2727 ( .I(addr_C1_M[14]), .ZN(n2417) );
  LVT_CLKNHSV0 U2728 ( .I(stateP2[1]), .ZN(n2465) );
  LVT_CLKNHSV0 U2729 ( .I(addr_C2_M[14]), .ZN(n2449) );
  LVT_CLKNHSV0 U2730 ( .I(addr_C1_M[0]), .ZN(n2415) );
  LVT_CLKNHSV0 U2731 ( .I(addr_P1_C1[0]), .ZN(n3059) );
  LVT_CLKNHSV0 U2732 ( .I(addr_C2_C1[13]), .ZN(n2412) );
  LVT_CLKNHSV0 U2733 ( .I(addr_C2_C1[14]), .ZN(n2403) );
  LVT_CLKNHSV0 U2734 ( .I(addr_C2_C1[5]), .ZN(n2466) );
  LVT_CLKNHSV0 U2735 ( .I(addr_C2_C1[9]), .ZN(n2467) );
  LVT_CLKNHSV0 U2736 ( .I(allowReadAddr_C2_C1[8]), .ZN(n2468) );
  LVT_CLKNHSV0 U2737 ( .I(allowReadAddr_C2_C1[7]), .ZN(n2469) );
  LVT_CLKNHSV0 U2738 ( .I(addr_C2_C1[12]), .ZN(n2560) );
  LVT_CLKNHSV0 U2739 ( .I(en_C2_P2), .ZN(n2464) );
  LVT_CLKNHSV0 U2740 ( .I(addr_C2_M[11]), .ZN(n2446) );
  LVT_CLKNHSV0 U2741 ( .I(addr_C2_M[13]), .ZN(n2445) );
  LVT_CLKNHSV0 U2742 ( .I(addr_C2_C1[6]), .ZN(n2559) );
  LVT_CLKNHSV1 U2743 ( .I(addr_C2_C1[7]), .ZN(n2558) );
  LVT_CLKNHSV0 U2744 ( .I(addr_C2_C1[11]), .ZN(n2556) );
  LVT_CLKNHSV0 U2745 ( .I(allowReadAddr_C2_C1[11]), .ZN(n2472) );
  LVT_CLKNHSV0 U2746 ( .I(addr_C2_M[4]), .ZN(n2444) );
  LVT_CLKNHSV0 U2747 ( .I(mb_stall), .ZN(n2474) );
  LVT_CLKNHSV0 U2748 ( .I(allowReadAddr_C2_C1[3]), .ZN(n2477) );
  LVT_CLKNHSV1 U2749 ( .I(allowReadAddr_C1_C2[6]), .ZN(n2481) );
  LVT_CLKNHSV0 U2750 ( .I(allowReadAddr_C2_C1[0]), .ZN(n2495) );
  LVT_CLKNHSV0 U2751 ( .I(addr_C2_M[7]), .ZN(n2442) );
  LVT_CLKNHSV0 U2752 ( .I(allowReadAddr_C2_C1[5]), .ZN(n2494) );
  LVT_CLKNHSV1 U2753 ( .I(addr_P1_C1[6]), .ZN(n2557) );
  LVT_CLKNHSV1 U2754 ( .I(allowReadAddr_C1_C2[7]), .ZN(n2471) );
  LVT_CLKNHSV0 U2755 ( .I(allowReadAddr_C2_C1[1]), .ZN(n2493) );
  LVT_CLKNHSV0 U2756 ( .I(allowReadAddr_C2_C1[2]), .ZN(n2492) );
  LVT_CLKNHSV0 U2757 ( .I(allowReadAddr_C2_C1[9]), .ZN(n2489) );
  LVT_CLKNHSV1 U2758 ( .I(allowReadAddr_C1_C2[14]), .ZN(n2475) );
  LVT_CLKNHSV1 U2759 ( .I(addr_P1_C1[13]), .ZN(n2575) );
  LVT_CLKNHSV1 U2760 ( .I(addr_P1_C1[7]), .ZN(n2514) );
  LVT_CLKNHSV1 U2761 ( .I(allowReadAddr_C1_C2[8]), .ZN(n2470) );
  LVT_CLKNHSV0 U2762 ( .I(allowReadAddr_C1_C2[0]), .ZN(n2500) );
  LVT_CLKNHSV0 U2763 ( .I(allowReadAddr_C2_C1[10]), .ZN(n2488) );
  LVT_CLKNHSV1 U2764 ( .I(addr_P1_C1[8]), .ZN(n2530) );
  LVT_CLKNHSV1 U2765 ( .I(allowReadAddr_C1_C2[13]), .ZN(n2476) );
  LVT_CLKNHSV0 U2766 ( .I(allowReadAddr_C2_C1[12]), .ZN(n2499) );
  LVT_CLKNHSV0 U2767 ( .I(addr_P1_C1[12]), .ZN(n2574) );
  LVT_CLKNHSV0 U2768 ( .I(allowReadAddr_C1_C2[9]), .ZN(n2491) );
  LVT_CLKNHSV0 U2769 ( .I(allowReadAddr_C1_C2[12]), .ZN(n2487) );
  LVT_CLKNHSV1 U2770 ( .I(addr_P1_C1[11]), .ZN(n2576) );
  LVT_CLKNHSV1 U2771 ( .I(allowReadAddr_C1_C2[11]), .ZN(n2473) );
  LVT_CLKNHSV1 U2772 ( .I(addr_P1_C1[9]), .ZN(n2531) );
  LVT_CLKNHSV0 U2773 ( .I(allowReadAddr_C1_C2[10]), .ZN(n2490) );
  LVT_CLKNHSV1 U2774 ( .I(addr_P1_C1[10]), .ZN(n2529) );
  LVT_CLKNHSV0 U2775 ( .I(addr_P1_C1[5]), .ZN(n2550) );
  LVT_CLKNHSV1 U2776 ( .I(addr_P1_C1[4]), .ZN(n2578) );
  LVT_CLKNHSV0 U2777 ( .I(allowReadAddr_C1_C2[5]), .ZN(n2496) );
  LVT_NOR2HSV0 U2778 ( .A1(ins_code2_proc2[22]), .A2(n2587), .ZN(n2583) );
  LVT_NOR2HSV0 U2779 ( .A1(ins_code1_proc1[22]), .A2(n2592), .ZN(n2589) );
  LVT_NOR2HSV2 U2780 ( .A1(n1674), .A2(n2950), .ZN(n2951) );
  LVT_BUFHSV2 U2781 ( .I(n2951), .Z(n3030) );
  LVT_BUFHSV2 U2782 ( .I(n2951), .Z(n3031) );
  LVT_INHSV2 U2783 ( .I(n2952), .ZN(n3028) );
  LVT_NOR2HSV2 U2784 ( .A1(n534), .A2(C2_stall), .ZN(n3001) );
  LVT_NAND2HSV0 U2785 ( .A1(n3015), .A2(n3001), .ZN(n2954) );
  LVT_NOR2HSV2 U2786 ( .A1(n2975), .A2(n2999), .ZN(n2984) );
  LVT_INHSV2 U2787 ( .I(n431), .ZN(n2389) );
  LVT_NOR2HSV2 U2788 ( .A1(n2984), .A2(n2389), .ZN(n3017) );
  LVT_INHSV2 U2789 ( .I(n3018), .ZN(n3022) );
  HVT_NAND3HSV0 U2790 ( .A1(n3022), .A2(n3023), .A3(n2955), .ZN(n1817) );
  LVT_INHSV2 U2791 ( .I(C1_addr_9_), .ZN(n2521) );
  LVT_INHSV2 U2792 ( .I(C1_addr_10_), .ZN(n2524) );
  LVT_INHSV2 U2793 ( .I(C1_addr_6_), .ZN(n2538) );
  LVT_INHSV2 U2794 ( .I(C1_addr_8_), .ZN(n2541) );
  LVT_INHSV2 U2795 ( .I(C1_addr_4_), .ZN(n2579) );
  LVT_INHSV2 U2796 ( .I(C1_addr_0_), .ZN(n3057) );
  LVT_INHSV2 U2797 ( .I(C1_addr_15_), .ZN(n2580) );
  LVT_INHSV2 U2798 ( .I(C1_addr_3_), .ZN(n2540) );
  LVT_INHSV2 U2799 ( .I(C1_addr_2_), .ZN(n2539) );
  LVT_INHSV2 U2800 ( .I(C1_addr_5_), .ZN(n2542) );
  LVT_INHSV2 U2801 ( .I(C1_addr_7_), .ZN(n2522) );
  LVT_INHSV2 U2802 ( .I(C1_addr_14_), .ZN(n2545) );
  LVT_INHSV2 U2803 ( .I(C1_addr_1_), .ZN(n2555) );
  LVT_INHSV2 U2804 ( .I(mb_chipSelect), .ZN(n2463) );
  LVT_INHSV2 U2805 ( .I(C2_addr_5_), .ZN(n2523) );
  LVT_INHSV2 U2806 ( .I(C2_addr_8_), .ZN(n3080) );
  LVT_INHSV2 U2807 ( .I(C2_addr_9_), .ZN(n2515) );
  LVT_INHSV2 U2808 ( .I(C2_addr_10_), .ZN(n2516) );
  LVT_INHSV2 U2809 ( .I(C2_addr_2_), .ZN(n2564) );
  LVT_INHSV2 U2810 ( .I(C2_addr_12_), .ZN(n2532) );
  LVT_INHSV2 U2811 ( .I(C2_addr_15_), .ZN(n2534) );
  LVT_INHSV2 U2812 ( .I(addr_P2_C2[8]), .ZN(n3088) );
  LVT_INHSV2 U2813 ( .I(addr_P2_C2[2]), .ZN(n3095) );
  LVT_INHSV2 U2814 ( .I(addr_P2_C2[1]), .ZN(n3089) );
  LVT_INHSV2 U2815 ( .I(addr_P2_C2[15]), .ZN(n3085) );
  LVT_INHSV2 U2816 ( .I(C2_addr_13_), .ZN(n2533) );
  LVT_INHSV2 U2817 ( .I(C2_addr_4_), .ZN(n2546) );
  LVT_INHSV2 U2818 ( .I(addr_P2_C2[10]), .ZN(n3093) );
  LVT_INHSV2 U2819 ( .I(addr_P2_C2[12]), .ZN(n3091) );
  LVT_INHSV2 U2820 ( .I(addr_P2_C2[5]), .ZN(n3087) );
  LVT_INHSV2 U2821 ( .I(addr_P2_C2[9]), .ZN(n3094) );
  LVT_INHSV2 U2822 ( .I(C2_addr_11_), .ZN(n2563) );
  LVT_INHSV2 U2823 ( .I(C2_addr_14_), .ZN(n2535) );
  LVT_INHSV2 U2824 ( .I(C2_addr_7_), .ZN(n3079) );
  LVT_INHSV2 U2825 ( .I(C2_addr_0_), .ZN(n3082) );
  LVT_INHSV2 U2826 ( .I(C2_addr_6_), .ZN(n3081) );
  LVT_INHSV2 U2827 ( .I(addr_P2_C2[13]), .ZN(n2562) );
  LVT_INHSV2 U2828 ( .I(addr_P2_C2[14]), .ZN(n2395) );
  LVT_INHSV2 U2829 ( .I(addr_P2_C2[11]), .ZN(n3086) );
  LVT_INHSV2 U2830 ( .I(addr_P2_C2[7]), .ZN(n3090) );
  LVT_INHSV2 U2831 ( .I(addr_P2_C2[6]), .ZN(n3096) );
  LVT_INHSV2 U2832 ( .I(addr_P2_C2[4]), .ZN(n3097) );
  LVT_NAND2HSV2 U2833 ( .A1(n591), .A2(n2957), .ZN(n1635) );
  LVT_AND2HSV2 U2834 ( .A1(n2958), .A2(n3067), .Z(n2988) );
  LVT_AND2HSV2 U2835 ( .A1(n2959), .A2(n2988), .Z(n2979) );
  LVT_NAND2HSV2 U2836 ( .A1(n2979), .A2(n3068), .ZN(n683) );
  LVT_INHSV2 U2837 ( .I(n683), .ZN(n3051) );
  LVT_NAND2HSV2 U2838 ( .A1(n534), .A2(n693), .ZN(n441) );
  LVT_CLKNHSV0 U2839 ( .I(n3065), .ZN(n2995) );
  LVT_AOI21HSV2 U2840 ( .A1(n2960), .A2(n2995), .B(n2969), .ZN(n2961) );
  LVT_OAI21HSV0 U2841 ( .A1(n2961), .A2(n641), .B(n3068), .ZN(n2962) );
  LVT_NAND2HSV2 U2842 ( .A1(n2962), .A2(n683), .ZN(n1560) );
  LVT_NAND2HSV2 U2843 ( .A1(n592), .A2(n2963), .ZN(n1662) );
  LVT_NAND2HSV2 U2844 ( .A1(n1662), .A2(n3068), .ZN(n2973) );
  LVT_NAND3HSV2 U2845 ( .A1(n2973), .A2(n683), .A3(n2964), .ZN(n1228) );
  LVT_CLKNAND2HSV1 U2846 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  LVT_NOR3HSV2 U2847 ( .A1(n2968), .A2(n1228), .A3(n2967), .ZN(n3048) );
  LVT_INHSV2 U2848 ( .I(n3048), .ZN(n1707) );
  LVT_INHSV2 U2849 ( .I(debugDelay[4]), .ZN(n2434) );
  LVT_INHSV2 U2850 ( .I(debugDelay[3]), .ZN(n2485) );
  LVT_NAND3HSV2 U2851 ( .A1(n2434), .A2(n2485), .A3(n2451), .ZN(n1451) );
  LVT_INHSV2 U2852 ( .I(n1451), .ZN(n2435) );
  LVT_INHSV2 U2853 ( .I(debugDelay[6]), .ZN(n2484) );
  LVT_INHSV2 U2854 ( .I(debugDelay[5]), .ZN(n2501) );
  LVT_NAND3HSV2 U2855 ( .A1(n2435), .A2(n2484), .A3(n2501), .ZN(n1434) );
  LVT_OAI21HSV2 U2856 ( .A1(n1662), .A2(n2969), .B(n3068), .ZN(n1664) );
  LVT_NAND3HSV2 U2857 ( .A1(n2979), .A2(n3055), .A3(rw_P1_C1[0]), .ZN(n2994)
         );
  LVT_INHSV2 U2858 ( .I(n2994), .ZN(n3040) );
  LVT_INHSV2 U2859 ( .I(n1228), .ZN(n3050) );
  LVT_NAND2HSV2 U2860 ( .A1(stateP1[0]), .A2(stateP1[1]), .ZN(n673) );
  LVT_NAND2HSV2 U2861 ( .A1(stateP2[1]), .A2(stateP2[0]), .ZN(n571) );
  LVT_NAND4HSV2 U2862 ( .A1(n3048), .A2(n2972), .A3(n2971), .A4(n2970), .ZN(
        n1569) );
  LVT_OAI21HSV2 U2863 ( .A1(n683), .A2(n3066), .B(n2973), .ZN(n1250) );
  LVT_INAND2HSV2 U2864 ( .A1(rw_P2_C2[1]), .B1(n3099), .ZN(n2974) );
  LVT_INAND3HSV2 U2865 ( .A1(n3073), .B1(n2975), .B2(n2974), .ZN(n3009) );
  LVT_OAI21HSV0 U2866 ( .A1(rw_C2_M[1]), .A2(n2452), .B(rw_C1_M[0]), .ZN(n2976) );
  LVT_IOA21HSV2 U2867 ( .A1(n707), .A2(rw_C2_M[0]), .B(n2976), .ZN(n1592) );
  LVT_IAO21HSV2 U2868 ( .A1(n2977), .A2(pc_proc2_code2[2]), .B(n2993), .ZN(
        P2_N106) );
  LVT_IAO21HSV2 U2869 ( .A1(n2978), .A2(pc_proc1_code1[2]), .B(n2991), .ZN(
        P1_N106) );
  LVT_INAND3HSV2 U2870 ( .A1(rw_P2_C2[1]), .B1(rw_P2_C2[0]), .B2(n3099), .ZN(
        n3024) );
  LVT_INOR2HSV1 U2871 ( .A1(n3024), .B1(n2394), .ZN(n449) );
  LVT_AND2HSV2 U2872 ( .A1(n2979), .A2(n3066), .Z(n2411) );
  LVT_INHSV2 U2873 ( .I(n3078), .ZN(n2986) );
  LVT_OAI211HSV0 U2874 ( .A1(n2982), .A2(n2981), .B(n2980), .C(n3098), .ZN(
        n2983) );
  LVT_OAI21HSV0 U2875 ( .A1(n3024), .A2(n3015), .B(n2983), .ZN(n2985) );
  LVT_AOI211HSV1 U2876 ( .A1(n3070), .A2(n2986), .B(n2985), .C(n2984), .ZN(
        n529) );
  LVT_OA31HSV2 U2877 ( .A1(n2989), .A2(n2988), .A3(n591), .B(n2987), .Z(n1655)
         );
  LVT_OA21HSV2 U2878 ( .A1(n2991), .A2(pc_proc1_code1[3]), .B(n2990), .Z(
        P1_N107) );
  LVT_OA21HSV2 U2879 ( .A1(n2993), .A2(pc_proc2_code2[3]), .B(n2992), .Z(
        P2_N107) );
  LVT_CLKNHSV0 U2880 ( .I(n2512), .ZN(n2996) );
  LVT_OAI211HSV1 U2881 ( .A1(n2996), .A2(n2995), .B(n683), .C(n2994), .ZN(n681) );
  LVT_CLKNHSV0 U2882 ( .I(n3015), .ZN(n2998) );
  LVT_OAI22HSV1 U2883 ( .A1(n3000), .A2(n2999), .B1(n2998), .B2(n2997), .ZN(
        n3002) );
  LVT_CLKNAND2HSV1 U2884 ( .A1(n3002), .A2(n3001), .ZN(n3016) );
  LVT_INAND2HSV0 U2885 ( .A1(n3003), .B1(n3070), .ZN(n3007) );
  LVT_AND2HSV2 U2886 ( .A1(n3016), .A2(n3007), .Z(n542) );
  HVT_OAI21HSV0 U2887 ( .A1(n3084), .A2(n1898), .B(n3004), .ZN(n3005) );
  LVT_NAND3HSV0 U2888 ( .A1(n3007), .A2(n3006), .A3(n3005), .ZN(n3008) );
  LVT_AOI211HSV1 U2889 ( .A1(msg_C2_C1), .A2(n3047), .B(n3008), .C(n3009), 
        .ZN(n495) );
  LVT_INHSV2 U2890 ( .I(n3009), .ZN(n3021) );
  LVT_NAND2HSV0 U2891 ( .A1(n3072), .A2(n3099), .ZN(n3010) );
  LVT_OAI211HSV1 U2892 ( .A1(n693), .A2(n694), .B(n3021), .C(n3010), .ZN(n501)
         );
  LVT_OA21HSV2 U2893 ( .A1(n3012), .A2(pc_proc1_code1[6]), .B(n3011), .Z(
        P1_N110) );
  LVT_OA21HSV2 U2894 ( .A1(n3014), .A2(pc_proc2_code2[6]), .B(n3013), .Z(
        P2_N110) );
  LVT_NAND2HSV2 U2895 ( .A1(n3073), .A2(n3015), .ZN(n3026) );
  LVT_INAND4HSV1 U2896 ( .A1(n536), .B1(n3026), .B2(n3017), .B3(n3016), .ZN(
        n425) );
  LVT_INHSV2 U2897 ( .I(n3023), .ZN(n3019) );
  LVT_AOI211HSV1 U2898 ( .A1(n3077), .A2(n3019), .B(n3018), .C(n440), .ZN(n692) );
  LVT_CLKNAND2HSV0 U2899 ( .A1(n440), .A2(n3070), .ZN(n3020) );
  LVT_OAI211HSV1 U2900 ( .A1(n3076), .A2(n417), .B(n3021), .C(n3020), .ZN(n442) );
  LVT_AND3HSV2 U2901 ( .A1(n3078), .A2(n3077), .A3(n3076), .Z(n3034) );
  LVT_INAND2HSV2 U2902 ( .A1(n441), .B1(n3027), .ZN(n732) );
endmodule

